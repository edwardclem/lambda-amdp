�� sr -edu.cornell.cs.nlp.spf.parser.ccg.model.Model�5B��B�~ L featureSetst Ljava/util/List;L independentLexicalFeatureSetsq ~ L invalidFeaturest Ljava/util/Set;L lexicont -Ledu/cornell/cs/nlp/spf/ccg/lexicon/ILexicon;L thetat 4Ledu/cornell/cs/nlp/spf/base/hashvector/IHashVector;xpsr &java.util.Collections$UnmodifiableList�%1�� L listq ~ xr ,java.util.Collections$UnmodifiableCollectionB ��^� L ct Ljava/util/Collection;xpsr java.util.LinkedList)S]J`�"  xpw   sr Pedu.cornell.cs.nlp.spf.parser.ccg.factoredlex.features.FactoredLexicalFeatureSet�g�պ��� D 
entryScaleI lexemeNextIdD lexemeScaleI nonFactoredNextIdI templateNextIdD templateScaleL entryInitialScorert :Ledu/cornell/cs/nlp/utils/collections/ISerializableScorer;L 	lexemeIdst 5Lit/unimi/dsi/fastutil/objects/Object2IntOpenHashMap;L lexemeInitialScorerq ~ L nonFactoredIdsq ~ L templateIdsq ~ L templateInitialScorerq ~ xr Iedu.cornell.cs.nlp.spf.parser.ccg.model.lexical.AbstractLexicalFeatureSetZ���n3�� Z computeSyntaxAttributeFeaturesL 
featureTagt Ljava/lang/String;L ignoreFiltert Ljava/util/function/Predicate;xp t FACLEXsr !java.lang.invoke.SerializedLambdaoaД,)6� 
I implMethodKind[ capturedArgst [Ljava/lang/Object;L capturingClasst Ljava/lang/Class;L functionalInterfaceClassq ~ L functionalInterfaceMethodNameq ~ L "functionalInterfaceMethodSignatureq ~ L 	implClassq ~ L implMethodNameq ~ L implMethodSignatureq ~ L instantiatedMethodTypeq ~ xp   ur [Ljava.lang.Object;��X�s)l  xp    vr 0edu.cornell.cs.nlp.utils.function.PredicateUtils           xpt java/util/function/Predicatet testt (Ljava/lang/Object;)Zt 0edu/cornell/cs/nlp/utils/function/PredicateUtilst lambda$alwaysTrue$bcad8f2c$1q ~ q ~ ?�         X?�             ?�������sr Eedu.cornell.cs.nlp.spf.parser.ccg.features.basic.scorer.UniformScorerQ�B���S D scorexp        sr 3it.unimi.dsi.fastutil.objects.Object2IntOpenHashMap         F fI sizexr 3it.unimi.dsi.fastutil.objects.AbstractObject2IntMap�o��K<z  xr 8it.unimi.dsi.fastutil.objects.AbstractObject2IntFunction�o��K<z I defRetValuexp    ?@     Xsr 9edu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.Lexeme	I����� I hashCodeCacheL 
attributesq ~ L 	constantsq ~ L 
propertiest Ljava/util/Map;L 	signaturet GLedu/cornell/cs/nlp/spf/ccg/lexicon/factored/lambda/FactoringSignature;L tokenst ,Ledu/cornell/cs/nlp/spf/base/token/TokenSeq;xp ��sr java.util.Collections$EmptyListz��<���  xpsq ~ q ~ -q ~ -sr %java.util.Collections$UnmodifiableMap��t�B L mq ~ (xpsq ~ /sr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t origint genlexxsr Eedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoringSignature�ڝ�U鞉 I hashCodeI numAttributesL typesq ~ xp  �    sq ~ sr java.util.ArrayListx����a� I sizexp    w    xq ~ :sr *edu.cornell.cs.nlp.spf.base.token.TokenSeq�py��An I hashCode[ tokenst [Ljava/lang/String;xp H�ur [Ljava.lang.String;��V��{G  xp   t Thew   Bsq ~ '~��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sr 0edu.cornell.cs.nlp.spf.mr.lambda.LogicalConstant=Q��� L baseNameq ~ L nameq ~ xr %edu.cornell.cs.nlp.spf.mr.lambda.Term�(G^� L typet .Ledu/cornell/cs/nlp/spf/mr/language/type/Type;xr 2edu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression
n�tL�h  xpsr 3edu.cornell.cs.nlp.spf.mr.language.type.ComplexType� �g��V L domainq ~ HL rangeq ~ Hxr ,edu.cornell.cs.nlp.spf.mr.language.type.Typeg���� I hashCodeCacheL nameq ~ xpgA�t <<e,t>,<<e,n>,e>>sq ~ K|-t <e,t>sr 0edu.cornell.cs.nlp.spf.mr.language.type.TermType��6��ǭ L parentt 2Ledu/cornell/cs/nlp/spf/mr/language/type/TermType;xq ~ L   et epsq ~ Q   tt tpsq ~ KH��t 	<<e,n>,e>sq ~ K|st <e,n>q ~ Ssq ~ Q   nt nq ~ Sq ~ St argmaxt argmax:<<e,t>,<<e,n>,e>>sq ~ Fq ~ Yt sizet 
size:<e,n>xq ~ Eq ~ Dsq ~ /sq ~ /sq ~ 2?@     w      q ~ 4t fixed_domainxsq ~ 6�C�j    sq ~ sq ~ 9   w   sq ~ KW�i�t <<e,t>,<<e,e>,e>>q ~ Osq ~ KHgKt 	<<e,e>,e>sq ~ K|\t <e,e>q ~ Sq ~ Sq ~ Sq ~ mxq ~ hsq ~ ;��uq ~ >   t largestw   %sq ~ '��q ~ -sq ~ sq ~ sq ~ 9   w   sq ~ Fsq ~ K?z��t 	<e,<e,n>>q ~ Sq ~ Yt distt dist:<e,<e,n>>xq ~ uq ~ tsq ~ /q ~ 1sq ~ 6?zy�    sq ~ sq ~ 9   w   sq ~ K?zu�t 	<e,<e,e>>q ~ Sq ~ mxq ~ ~sq ~ ; /#�uq ~ >   t doorw   Msq ~ ' 3�Nq ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~ �sq ~ ; 3<uq ~ >   t movew   Dsq ~ '�FĘsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ Fsq ~ K?z�t 	<e,<e,t>>q ~ Sq ~ Ot int in:<e,<e,t>>xq ~ �q ~ �sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~ �sq ~ ;  cuq ~ >   q ~ �w   sq ~ 'X�7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ Fq ~ Mt argmint argmin:<<e,t>,<<e,n>,e>>q ~ vxq ~ �q ~ �sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6�BQ�    sq ~ sq ~ 9   w   q ~ iq ~ xq ~ �sq ~ ;A#�"uq ~ >   t closestt tow   sq ~ '�lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �q ~ _xq ~ �q ~ �sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6�C�j    sq ~ sq ~ 9   w   q ~ iq ~ mxq ~ �sq ~ ;��]uq ~ >   t smallestw   !sq ~ '}g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ Fq ~ Ot agentt agent:<e,t>xq ~ �q ~ �sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~ �sq ~ ;�CCuq ~ >   q ~ �w   sq ~ 'w���q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~ �q ~ �sq ~ /q ~ 1sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~ �sq ~ ; zuq ~ >   t andw   Ssq ~ '�kgdq ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~ �q ~ �sq ~ /q ~ 1sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~ �sq ~ ; $�/uq ~ >   t Movew   4sq ~ '�b�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ Fq ~ Ot blockt block:<e,t>xq ~ �q ~ �sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~ �sq ~ ;���uq ~ >   q ~ �w   sq ~ 'l�8q ~ -sq ~ sq ~ sq ~ 9   w   sq ~ Fq ~ Ot greent green:<e,t>xq ~ �q ~ �sq ~ /q ~ 1sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~ �sq ~ ;��Auq ~ >   q ~ �w   2sq ~ '�b�q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ �xq ~q ~sq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~	sq ~ ;  	Fuq ~ >   t Gow   .sq ~ ';��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ Fq ~ Ot roomt 
room:<e,t>xq ~q ~sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~sq ~ ; 5�uq ~ >   q ~w   
sq ~ '�CZ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �q ~ �xq ~!q ~ sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6�C�;    sq ~ sq ~ 9   w   q ~ iq ~ Oxq ~'sq ~ ;l�0�uq ~ >   t nearestw   'sq ~ '  ��q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~0sq ~ ;  �uq ~ >   q ~ �w   1sq ~ 'w�(sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~7q ~6sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~=sq ~ ; �suq ~ >   t goq ~ �w   sq ~ ' �|q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~Fsq ~ ; \=uq ~ >   t Youw   6sq ~ '{k��q ~ Bsq ~ sq ~ sq ~ 
w   q ~ Jxq ~Mq ~Lsq ~ /q ~ csq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~Qq ~ ow   sq ~ 'C�;zq ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~Uq ~Tsq ~ /q ~#sq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~Yq ~(w   	sq ~ '�X�\q ~sq ~ sq ~ sq ~ 
w   q ~ vq ~ �xq ~]q ~\sq ~ /q ~#sq ~ 6�Pi�    sq ~ sq ~ 9   w   q ~ q ~ Oxq ~aq ~(w   sq ~ '�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �q ~ �xq ~fq ~esq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6�C�;    sq ~ sq ~ 9   w   q ~ iq ~ Oxq ~lsq ~ ;3�N�uq ~ >   q ~ �w   )sq ~ 'Es�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �q ~ vxq ~sq ~rsq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6�BQ�    sq ~ sq ~ 9   w   q ~ iq ~ xq ~ysq ~ ;-��uq ~ >   q ~*q ~ �w   sq ~ '��;q ~ �sq ~ sq ~ sq ~ 
w   q ~ �xq ~q ~~sq ~ /q ~ �sq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~�q ~ �w   sq ~ '�X�q ~ -sq ~ sq ~ sq ~ 9   w   sq ~ Fq ~ Oq ~ �t 
door:<e,t>xq ~�q ~�sq ~ /q ~ 1sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~�sq ~ ;l�0�uq ~ >   q ~*w   Jsq ~ 'ǋ�q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ �xq ~�q ~�sq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~�sq ~ ; )'uq ~ >   t Walkw   ;sq ~ ' �-q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ; �uq ~ >   t Canw   9sq ~ '�F��q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~�q ~�sq ~ /q ~ 1sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~�q ~1w   ,sq ~ '�{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~�sq ~ ;4P�uq ~ >   q ~ �q ~ �w   (sq ~ ' L�q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ; �]uq ~ >   t youw   :sq ~ '  ��q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ;  iuq ~ >   t itw   Usq ~ '�F�{q ~ -sq ~ q ~�q ~�sq ~ /q ~ 1sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~�q ~
w   0sq ~ 'y�M�q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ �xq ~�q ~�sq ~ /q ~ 1sq ~ 6�C�;    sq ~ sq ~ 9   w   q ~ iq ~ Oxq ~�q ~ �w   Lsq ~ '��q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ vxq ~�q ~�sq ~ /q ~ 1sq ~ 6�BQ�    sq ~ sq ~ 9   w   q ~ iq ~ xq ~�q ~ �w   Ksq ~ '���q ~ -sq ~ sq ~ sq ~ 9   w   sq ~ Fq ~ �t next_tot next_to:<e,<e,t>>xq ~�q ~�sq ~ /q ~ 1sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~�sq ~ ; 3�1uq ~ >   t nextw   Fsq ~ ' 0�nsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ; 0R/uq ~ >   t canq ~�w   sq ~ '��
q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~ q ~�sq ~ /q ~ 1sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~sq ~ ;�R�uq ~ >   t 
containingw   Gsq ~ 'H��q ~ �sq ~ sq ~ sq ~ 
w   q ~ _xq ~q ~
sq ~ /q ~ �sq ~ 6|!<    sq ~ sq ~ 9   w   q ~ mxq ~q ~ �w   $sq ~ ' 8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6  �    sq ~ sq ~ 9    w    xq ~sq ~ ; ��uq ~ >   t thew   sq ~ '�b�q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ �xq ~!q ~ sq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~%sq ~ ;  &uq ~ >   q ~@w   8sq ~ '���Lq ~csq ~ sq ~ sq ~ 
w   q ~ �xq ~+q ~*sq ~ /q ~hsq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~/q ~mw   sq ~ 'I�kq ~csq ~ sq ~ sq ~ 
w   q ~ vxq ~3q ~2sq ~ /q ~hsq ~ 6?zy�    sq ~ sq ~ 9   w   q ~ xq ~7q ~mw   sq ~ '䳙Qq ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~;q ~:sq ~ /q ~#sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~?q ~(w   sq ~ '��F;q ~sq ~ sq ~ sq ~ 
w   q ~ �q ~ vq ~ �xq ~Cq ~Bsq ~ /q ~#sq ~ 6���    sq ~ sq ~ 9   w   q ~ iq ~ q ~ Oxq ~Gq ~(w   sq ~ '�y�Dq ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~Kq ~Jsq ~ /q ~ 1sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~Osq ~ ; 3<uq ~ >   q ~ �w   Tsq ~ 'Ǔoq ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ �xq ~Uq ~Tsq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~Ysq ~ ; 1f�uq ~ >   t intow   Asq ~ '�Ҭq ~ -sq ~ sq ~ sq ~ 9   w   q ~ vq ~ �xq ~`q ~_sq ~ /q ~ 1sq ~ 6�Pi�    sq ~ sq ~ 9   w   q ~ q ~ Oxq ~dq ~ �w   Qsq ~ 'x��q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~hq ~gsq ~ /q ~ 1sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~lq ~ �w   Psq ~ '��6�q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ �xq ~pq ~osq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~tsq ~ ;�e.=uq ~ >   t yourselfw   >sq ~ '����q ~ -sq ~ sq ~ sq ~ 9   w   q ~�q ~ �xq ~{q ~zsq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~sq ~ ; 3�1uq ~ >   q ~�w   Esq ~ '�b8q ~ -sq ~ q ~q ~sq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~�q ~1w   +sq ~ '�HY�q ~4sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ /q ~9sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~�q ~>w   sq ~ '�@�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ;�@(uq ~ >   t pleasew   sq ~ ' +�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ; �Muq ~ >   t putw   sq ~ '��.�q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~�q ~�sq ~ /q ~ 1sq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~�q ~ �w   Osq ~ '~�_q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ /q ~�sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~�q ~�w   sq ~ 'ǆ��q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ �xq ~�q ~�sq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~�q ~ �w   3sq ~ 'WS�q ~ �sq ~ sq ~ sq ~ 
w   q ~ vxq ~�q ~�sq ~ /q ~ �sq ~ 6?zy�    sq ~ sq ~ 9   w   q ~ xq ~�q ~ �w   sq ~ 'w�wnq ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~�q ~�sq ~ /q ~ 1sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~�q ~1w   -sq ~ '�q�&q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~�q ~�sq ~ /q ~ 1sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~�sq ~ ;�+�uq ~ >   t shouldw   Csq ~ ' %(nq ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ; $�/uq ~ >   q ~ �w   =sq ~ ' �lq ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ; ;-uq ~ >   t Putw   5sq ~ '  ��q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�q ~
w   *sq ~ '�c��q ~4sq ~ sq ~ sq ~ 
w   q ~ �q ~ �xq ~�q ~�sq ~ /q ~9sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~�q ~>w    sq ~ '3���q ~ Bsq ~ sq ~ sq ~ 
w   q ~ _xq ~q ~ sq ~ /q ~ csq ~ 6|!<    sq ~ sq ~ 9   w   q ~ mxq ~q ~ ow   sq ~ 'J��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ Fq ~ Ot bluet 
blue:<e,t>xq ~
q ~	sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~sq ~ ; .0�uq ~ >   q ~w    sq ~ '�+�0q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~sq ~ ;�+�uq ~ >   q ~�w   7sq ~ ' 1��q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~#sq ~ ; 1f�uq ~ >   q ~\w   Vsq ~ 'O9�q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ vq ~ �xq ~)q ~(sq ~ /q ~ 1sq ~ 6���    sq ~ sq ~ 9   w   q ~ iq ~ q ~ Oxq ~-q ~ �w   Nsq ~ '͖Y)q ~�sq ~ sq ~ sq ~ 
w   q ~ �q ~ �xq ~1q ~0sq ~ /q ~�sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~5q ~�w   sq ~ ' "v�q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~;sq ~ ; !��uq ~ >   t Grabw   Wsq ~ ' ��q ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~Dsq ~ ; tuq ~ >   t Getw   Rsq ~ 'XΖxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ Fq ~ Ot redt 	red:<e,t>xq ~Lq ~Ksq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~Usq ~ ; ��uq ~ >   q ~Nw   sq ~ '��mq ~ -sq ~ sq ~ sq ~ 9   w   q ~ �xq ~[q ~Zsq ~ /q ~ 1sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~_sq ~ ;���8uq ~ >   t thatt containsw   Hsq ~ 'rK�q ~ -sq ~ sq ~ sq ~ 9   w   q ~�xq ~gq ~fsq ~ /q ~ 1sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~ksq ~ ; /#�uq ~ >   q ~ �w   @sq ~ 'R+�Wq ~csq ~ sq ~ sq ~ 
w   q ~ vq ~ �xq ~qq ~psq ~ /q ~hsq ~ 6�Pi�    sq ~ sq ~ 9   w   q ~ q ~ Oxq ~uq ~mw   "sq ~ 'ǖE�q ~ -sq ~ sq ~ sq ~ 9   w   q ~ �q ~ �xq ~yq ~xsq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~}sq ~ ; 4=uq ~ >   t overw   ?sq ~ 'U��q ~psq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ /q ~usq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~�q ~zw   sq ~ '�G��q ~sq ~ sq ~ sq ~ 
w   q ~ �q ~ vxq ~�q ~�sq ~ /q ~#sq ~ 6�BQ�    sq ~ sq ~ 9   w   q ~ iq ~ xq ~�q ~(w   #sq ~ 'KԬq ~csq ~ sq ~ sq ~ 
w   q ~ �q ~ vxq ~�q ~�sq ~ /q ~hsq ~ 6�BQ�    sq ~ sq ~ 9   w   q ~ iq ~ xq ~�q ~mw   sq ~ '���pq ~sq ~ sq ~ sq ~ 
w   q ~ vxq ~�q ~�sq ~ /q ~#sq ~ 6?zy�    sq ~ sq ~ 9   w   q ~ xq ~�q ~(w   sq ~ '� q ~ �sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ /q ~ �sq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~�q ~ �w   sq ~ 'Cw��q ~psq ~ sq ~ sq ~ 
w   q ~ vxq ~�q ~�sq ~ /q ~usq ~ 6?zy�    sq ~ sq ~ 9   w   q ~ xq ~�q ~zw   sq ~ '��d6q ~csq ~ sq ~ sq ~ 
w   q ~ �q ~ vq ~ �xq ~�q ~�sq ~ /q ~hsq ~ 6���    sq ~ sq ~ 9   w   q ~ iq ~ q ~ Oxq ~�q ~mw   &sq ~ '�qxq ~ -sq ~ q ~ -q ~ -sq ~ /q ~ 1sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~ ;��9uq ~ >   t Carryw   <sq ~ '
iYuq ~csq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ /q ~hsq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~�q ~mw   sq ~ '�~��q ~ -sq ~ sq ~ sq ~ 9   w   q ~�q ~ �xq ~�q ~�sq ~ /q ~ 1sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~�sq ~ ; )'uq ~ >   q ~�w   Isq ~ 'w�q�q ~ -sq ~ q ~�q ~�sq ~ /q ~ 1sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~�q ~
w   /xsq ~ !        sq ~ #    ?@      xsq ~ #    ?@     sr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.LexicalTemplateg��%��	 I hashCodeL 	argumentsq ~ L 
propertiesq ~ (L 	signatureq ~ )L templatet 0Ledu/cornell/cs/nlp/spf/ccg/categories/Category;xpIH�xsq ~ sq ~ sq ~ 
w   sq ~ Fq ~ Ot #0<e,t>t #0<e,t>:<e,t>xq ~�q ~�sq ~ /q ~sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~�sr 5edu.cornell.cs.nlp.spf.ccg.categories.ComplexCategory�f�Ք�nl I hashCodeCacheL syntaxt <Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/ComplexSyntax;xr .edu.cornell.cs.nlp.spf.ccg.categories.CategorycK=�.A� L 	semanticst Ljava/lang/Object;xpsr 'edu.cornell.cs.nlp.spf.mr.lambda.Lambda��Kβ�� L argumentt +Ledu/cornell/cs/nlp/spf/mr/lambda/Variable;L bodyt 4Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L typet 5Ledu/cornell/cs/nlp/spf/mr/language/type/ComplexType;xq ~ Isr )edu.cornell.cs.nlp.spf.mr.lambda.Variable�u#$rP L 	singletonq ~ xq ~ Gq ~ Osr 5it.unimi.dsi.fastutil.objects.ReferenceSets$Singleton�7y�J| L elementq ~�xpq ~�sq ~�sq ~�q ~ Ssq ~�q ~�sr (edu.cornell.cs.nlp.spf.mr.lambda.Literalŕtb��� [ 	argumentst 5[Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L 	predicateq ~�[ 	signaturet /[Ledu/cornell/cs/nlp/spf/mr/language/type/Type;L typeq ~ Hxq ~ Iur 5[Ledu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression;|�㰢�[i  xp   sq ~�uq ~�   q ~�q ~�q ~�ur /[Ledu.cornell.cs.nlp.spf.mr.language.type.Type;>L5��  xp   q ~ Sq ~ Usq ~�uq ~�   q ~�sr ;it.unimi.dsi.fastutil.objects.ReferenceSets$UnmodifiableSet�7y�J|  xr Iit.unimi.dsi.fastutil.objects.ReferenceCollections$UnmodifiableCollection�7y�J| L 
collectiont 3Lit/unimi/dsi/fastutil/objects/ReferenceCollection;xpsr 2it.unimi.dsi.fastutil.objects.ReferenceOpenHashSet         F fI sizexp?@     q ~�q ~�xq ~�uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~�q ~�xsq ~ Fsr <edu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType&��M
� I minArgsZ orderSensitiveL optiont ELedu/cornell/cs/nlp/spf/mr/language/type/RecursiveComplexType$Option;xq ~ Kl�6�t <t*,t>q ~ Uq ~ U    sr Cedu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType$Option�^g� �� Z isOrderSensitiveI 
minNumArgsxp    q ~ �t 
and:<t*,t>uq ~   q ~ Uq ~ Uq ~ Usq ~sq ~?@     q ~�xq ~ Osr 4it.unimi.dsi.fastutil.objects.ReferenceSets$EmptySet�7y�J|  xpsq ~ KJW`Lt <<e,t>,<e,t>>q ~ Oq ~ OR:L]sr :edu.cornell.cs.nlp.spf.ccg.categories.syntax.ComplexSyntax$���q\P^ I hashCodeI 	numSlahesL leftt 5Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax;L rightq ~ L slasht 4Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Slash;xr 3edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntaxʊ�	�|��  xp�z�M   sr @edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntax$SimpleSyntax��eBg� I hashCodeL 	attributeq ~ L labelq ~ xq ~" 3�kt nonet Nq ~%sr 2edu.cornell.cs.nlp.spf.ccg.categories.syntax.Slashѕ�����> C cxp /w   sq ~�/�sq ~ sq ~ sq ~ 
w   sq ~ Fq ~ it #0<<e,t>,<<e,e>,e>>t %#0<<e,t>,<<e,e>,e>>:<<e,t>,<<e,e>,e>>sq ~ Fq ~ t #0<e,<e,e>>t #0<e,<e,e>>:<e,<e,e>>xq ~-q ~,sq ~ /q ~#sq ~ 6�BQ�    sq ~ sq ~ 9   w   q ~ iq ~ xq ~7sq ~�sq ~�sq ~�q ~ Osq ~�q ~:sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~?sq ~�uq ~�   q ~?sq ~sq ~?@     q ~:q ~?xq ~:uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~:xq ~ Osq ~�sq ~�q ~ Ssq ~�q ~Isq ~�uq ~�   sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~Psq ~�uq ~�   q ~Pq ~Qq ~ �uq ~   q ~ Sq ~ Uq ~q ~ Oq ~sq ~ Fsq ~ KI:��t 	<<e,t>,e>q ~ Oq ~ Sq ~t the:<<e,t>,e>uq ~   q ~ Oq ~ Sq ~Iq ~Jq ~1uq ~   q ~ Sq ~ Sq ~ Sq ~q ~ mq ~Fq ~.uq ~   q ~ Oq ~ mq ~ Sq ~q ~V~p�Nsq ~�ƥ�   sq ~$ 4�wq ~&t NPq ~%sq ~( \w   sq ~����sq ~ sq ~ sq ~ 
w    xq ~cq ~bsq ~ /q ~�sq ~ 6  �    sq ~ sq ~ 9    w    xq ~gsq ~�sq ~�sq ~�q ~ Usq ~�q ~jq ~jq ~sq ~ K��t <t,t>q ~ Uq ~ U���sq ~�|��   sq ~$ 3�q ~&t Sq ~oq ~)w   sq ~��9gsq ~ sq ~ sq ~ 
w   q ~.xq ~tq ~ssq ~ /q ~usq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~xsq ~�sq ~�sq ~�q ~ Ssq ~�q ~{sq ~�sq ~�q ~ Osq ~�q ~~sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�sq ~sq ~?@     q ~~q ~�xq ~~uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~~xq ~ Osq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~{q ~�sq ~sq ~?@     q ~�q ~{xq ~ vuq ~   q ~ Sq ~ Sq ~ [sq ~sq ~?@     q ~{xq ~ Ysq ~sq ~?@     q ~~q ~{xq ~.uq ~   q ~ Oq ~ mq ~ Ssq ~sq ~?@     q ~{xq ~Vq ~sq ~ Ke5Et <e,<<e,t>,e>>q ~ Sq ~Vj���sq ~�   sq ~�ƥ�   q ~]q ~%q ~_q ~]q ~)w   sq ~�(W~sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ /q ~sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~�sq ~�sq ~�q ~ Osq ~�q ~�sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�sq ~sq ~?@     q ~�q ~�xq ~�uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~�xq ~ Oq ~q ~(S�sq ~�z�M   q ~%q ~%q ~)w   sq ~ݎ���sq ~ sq ~ sq ~ 
w   q ~.sq ~ Fq ~ mt #0<e,e>t #0<e,e>:<e,e>xq ~�q ~�sq ~ /q ~ �sq ~ 6�C�j    sq ~ sq ~ 9   w   q ~ iq ~ mxq ~�sq ~�sq ~�sq ~�q ~ Osq ~�q ~�sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�sq ~sq ~?@     q ~�q ~�xq ~�uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~�xq ~ Osq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�uq ~   q ~ Sq ~ Sq ~q ~ mq ~�q ~.uq ~   q ~ Oq ~ mq ~ Sq ~q ~VZ`O�sq ~�ƥY   q ~]q ~%q ~)w   sq ~�A["fsq ~ sq ~ sq ~ 
w   q ~.xq ~�q ~�sq ~ /q ~#sq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~�sq ~�sq ~�q ~:sq ~�uq ~�   q ~>sq ~�q ~Isq ~�uq ~�   q ~Mq ~Iq ~Jq ~ vuq ~   q ~ Sq ~ Sq ~ [q ~q ~ Yq ~Fq ~.uq ~   q ~ Oq ~ mq ~ Sq ~q ~V�ړ�q ~\w   	sq ~�ێ8Msq ~ sq ~ sq ~ 
w   q ~.xq ~�q ~�sq ~ /q ~ �sq ~ 6W�m�    sq ~ sq ~ 9   w   q ~ ixq ~�sq ~�sq ~�q ~�sq ~�uq ~�   q ~�sq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~ _uq ~   q ~ Sq ~ [q ~q ~ Yq ~�q ~.uq ~   q ~ Oq ~ mq ~ Sq ~q ~Vy��q ~�w   
sq ~��/�lsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ /q ~ csq ~ 6|!<    sq ~ sq ~ 9   w   q ~ mxq ~sq ~�sq ~�sq ~�q ~ Osq ~�q ~sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~
sq ~�uq ~�   q ~
sq ~sq ~?@     q ~
q ~xq ~uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~xq ~ Osq ~�sq ~�q ~ Ssq ~�q ~sq ~�uq ~�   q ~q ~q ~�uq ~   q ~ Sq ~ Sq ~q ~ mq ~q ~ Juq ~   q ~ Oq ~ Yq ~ Sq ~q ~V�+@sq ~�ƥY   q ~]q ~%q ~)w   sq ~�oU��sq ~ sq ~ sq ~ 
w   q ~.q ~1xq ~q ~sq ~ /q ~usq ~ 6�BQ�    sq ~ sq ~ 9   w   q ~ iq ~ xq ~"sq ~�sq ~�q ~{sq ~�q ~~sq ~�uq ~�   q ~�sq ~�q ~�sq ~�uq ~�   q ~{q ~�sq ~sq ~?@     q ~�q ~{xq ~1uq ~   q ~ Sq ~ Sq ~ Ssq ~sq ~?@     q ~{xq ~ msq ~sq ~?@     q ~~q ~{xq ~.uq ~   q ~ Oq ~ mq ~ Ssq ~sq ~?@     q ~{xq ~Vq ~q ~����q ~�w   sq ~�I�psq ~ sq ~ sq ~ 
w   sq ~ Fq ~ �t #0<e,<e,t>>t #0<e,<e,t>>:<e,<e,t>>xq ~8q ~7sq ~ /q ~ �sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~?sq ~�sq ~�sq ~�q ~ Ssq ~�q ~Bsq ~�sq ~�q ~ Ssq ~�q ~Esq ~�uq ~�   q ~Eq ~Bsq ~sq ~?@     q ~Bq ~Exq ~9uq ~   q ~ Sq ~ Sq ~ Usq ~sq ~?@     q ~Bxq ~ Oq ~q ~ �H�o�sq ~�P�   sq ~$ 4��q ~&t PPq ~]q ~)w   sq ~ݍ'��sq ~ sq ~ sq ~ 
w   q ~.q ~1q ~�xq ~Tq ~Ssq ~ /q ~#sq ~ 6���    sq ~ sq ~ 9   w   q ~ iq ~ q ~ Oxq ~Xsq ~�sq ~�q ~:sq ~�uq ~�   q ~>sq ~�q ~Isq ~�uq ~�   sq ~�uq ~�   sq ~�q ~Psq ~�uq ~�   q ~Pq ~Qq ~�uq ~   q ~ Sq ~ Uq ~q ~ Oq ~q ~Uuq ~   q ~ Oq ~ Sq ~Iq ~Jq ~1uq ~   q ~ Sq ~ Sq ~ Sq ~q ~ mq ~Fq ~.uq ~   q ~ Oq ~ mq ~ Sq ~q ~V���q ~\w   sq ~݌?kisq ~ sq ~ sq ~ 
w    xq ~lq ~ksq ~ /q ~�sq ~ 6  �    sq ~ sq ~ 9    w    xq ~psq ~�sq ~�sq ~�q ~ Ssq ~�q ~ssq ~�sq ~�q ~ Osq ~�q ~vsq ~�uq ~�   q ~ssq ~sq ~?@     q ~sq ~vxq ~vuq ~   q ~ Sq ~ Usq ~sq ~?@     q ~sxsq ~ KI:�et 	<<e,t>,t>q ~ Oq ~ Uq ~sq ~ Ke5}\t <e,<<e,t>,t>>q ~ Sq ~�?g�sq ~+���   sq ~ȡ>Z   q ~oq ~Oq ~)q ~]q ~)w   sq ~�(�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~�sq ~�sq ~�q ~ Osq ~�q ~�sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�sq ~sq ~?@     q ~�q ~�xq ~�uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~�xq ~ Oq ~q ~(�>sq ~�|��   q ~oq ~oq ~)w   sq ~�ܞD�sq ~ sq ~ sq ~ 
w   q ~1q ~�xq ~�q ~�sq ~ /q ~hsq ~ 6�Pi�    sq ~ sq ~ 9   w   q ~ q ~ Oxq ~�sq ~�sq ~�sq ~�q ~ Osq ~�q ~�sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�sq ~sq ~?@     q ~�q ~�xq ~�uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~�xq ~ Osq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�uq ~   q ~ Sq ~ Uq ~q ~ Oq ~q ~Uuq ~   q ~ Oq ~ Sq ~�q ~�q ~1uq ~   q ~ Sq ~ Sq ~ Sq ~q ~ mq ~�q ~ �uq ~   q ~ Oq ~ Yq ~ Sq ~q ~V-��Hsq ~�ƥ�   q ~]q ~%q ~_w   sq ~����sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ /q ~�sq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~�sq ~�sq ~�q ~ Usq ~�q ~�q ~�q ~q ~l���sq ~�|�   q ~oq ~oq ~_w   sq ~�x�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ /sq ~ /sq ~ 2?@     w      q ~ 4q ~ exsq ~ 6  �    sq ~ sq ~ 9    w    xq ~�sq ~�sq ~�sq ~�q ~ Osq ~�q ~�sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�sq ~sq ~?@     q ~�q ~�xq ~�uq ~   q ~ Sq ~ Usq ~sq ~?@     q ~�xq ~ Oq ~�q ~Uuq ~   q ~ Oq ~ Sq ~q ~Vx~'sq ~�ƥY   q ~]q ~%q ~)w   sq ~�VN:�sq ~ sq ~ sq ~ 
w   q ~1xq ~�q ~�sq ~ /q ~hsq ~ 6?zy�    sq ~ sq ~ 9   w   q ~ xq ~�sq ~�sq ~�q ~�sq ~�uq ~�   q ~�sq ~�q ~�sq ~�uq ~�   sq ~�uq ~�   sq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~ �uq ~   q ~ Sq ~ Uq ~q ~ Oq ~q ~Uuq ~   q ~ Oq ~ Sq ~�q ~�q ~1uq ~   q ~ Sq ~ Sq ~ Sq ~q ~ mq ~�q ~ �uq ~   q ~ Oq ~ Yq ~ Sq ~q ~V�o��q ~�w   sq ~�^�>sq ~ sq ~ sq ~ 
w   q ~.q ~�xq ~q ~
sq ~ /q ~#sq ~ 6�C�;    sq ~ sq ~ 9   w   q ~ iq ~ Oxq ~sq ~�sq ~�q ~:sq ~�uq ~�   q ~>sq ~�q ~Isq ~�uq ~�   sq ~�uq ~�   sq ~�q ~Psq ~�uq ~�   q ~Pq ~Qq ~�uq ~   q ~ Sq ~ Uq ~q ~ Oq ~q ~Uuq ~   q ~ Oq ~ Sq ~Iq ~Jq ~ vuq ~   q ~ Sq ~ Sq ~ [q ~q ~ Yq ~Fq ~.uq ~   q ~ Oq ~ mq ~ Sq ~q ~Vz�Wq ~\w   sq ~��*z5sq ~ sq ~ sq ~ 
w   q ~9q ~�xq ~#q ~"sq ~ /q ~9sq ~ 6�W;    sq ~ sq ~ 9   w   q ~ �q ~ Oxq ~'sq ~�sq ~�sq ~�q ~ Ssq ~�q ~*sq ~�uq ~�   sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~1sq ~�uq ~�   q ~1q ~2q ~�uq ~   q ~ Sq ~ Uq ~q ~ Oq ~q ~Uuq ~   q ~ Oq ~ Sq ~*q ~+q ~9uq ~   q ~ Sq ~ Sq ~ Uq ~q ~ O���.sq ~ȠU�   q ~oq ~]q ~)w   sq ~݅*�sq ~ sq ~ sq ~ 
w   q ~�xq ~<q ~;sq ~ /q ~hsq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~@sq ~�sq ~�q ~�sq ~�uq ~�   q ~�sq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�q ~ vuq ~   q ~ Sq ~ Sq ~ [q ~q ~ Yq ~�q ~ �uq ~   q ~ Oq ~ Yq ~ Sq ~q ~V���q ~�w    sq ~���sq ~ sq ~ sq ~ 
w   q ~1xq ~Mq ~Lsq ~ /q ~ �sq ~ 6?zy�    sq ~ sq ~ 9   w   q ~ xq ~Qsq ~�sq ~�sq ~�q ~ Ssq ~�q ~Tsq ~�sq ~�q ~ Osq ~�q ~Wsq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~\sq ~�uq ~�   q ~\sq ~sq ~?@     q ~Wq ~\xq ~Wuq ~   q ~ Sq ~ Usq ~sq ~?@     q ~Wxq ~ Osq ~�sq ~�q ~ Ssq ~�q ~fsq ~�uq ~�   q ~Tq ~fsq ~sq ~?@     q ~Tq ~fxq ~1uq ~   q ~ Sq ~ Sq ~ Ssq ~sq ~?@     q ~Txq ~ msq ~sq ~?@     q ~Wq ~Txq ~ �uq ~   q ~ Oq ~ Yq ~ Ssq ~sq ~?@     q ~Txq ~Vq ~q ~�)�Xsq ~�   sq ~�ƥ�   q ~]q ~%q ~_q ~]q ~)w   sq ~�t�,sq ~ sq ~ sq ~ 
w   q ~9xq ~yq ~xsq ~ /q ~9sq ~ 6?z��    sq ~ sq ~ 9   w   q ~ �xq ~}sq ~�sq ~�q ~*sq ~�uq ~�   sq ~�uq ~�   sq ~�q ~1sq ~�uq ~�   q ~1q ~2q ~ �uq ~   q ~ Sq ~ Uq ~q ~ Oq ~q ~Uuq ~   q ~ Oq ~ Sq ~*q ~+q ~9uq ~   q ~ Sq ~ Sq ~ Uq ~q ~ Ot��q ~8w   sq ~ݵdZsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ /q ~ �sq ~ 6|!<    sq ~ sq ~ 9   w   q ~ mxq ~�sq ~�sq ~�q ~�sq ~�uq ~�   q ~�sq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�uq ~   q ~ Sq ~ Sq ~q ~ mq ~�q ~ �uq ~   q ~ Oq ~ Yq ~ Sq ~q ~Vn_E.q ~�w   sq ~���'sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ /q ~ �sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~�sr 4edu.cornell.cs.nlp.spf.ccg.categories.SimpleCategory��4_C� I hashCodeCacheL syntaxt BLedu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax$SimpleSyntax;xq ~�sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�uq ~   q ~ Sq ~ Uq ~q ~ O�Ǵq ~%w   sq ~��7�'sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ /q ~�sq ~ 6|#    sq ~ sq ~ 9   w   q ~ Oxq ~�sq ~�sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   sq ~�uq ~�   sq ~�sq ~�q ~ Ssq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�uq ~   q ~ Sq ~ Uq ~q ~ Oq ~q ~Uuq ~   q ~ Oq ~ Sq ~�q ~�q ~ �uq ~   q ~ Sq ~ Sq ~ Uq ~q ~ O�).sq ~ȠU�   q ~oq ~]q ~)w   xsq ~ !        sr Yedu.cornell.cs.nlp.spf.parser.ccg.features.lambda.LogicalExpressionCoordinationFeatureSet�4tHWcg+ Z cpapFeaturesZ cpp1FeaturesZ reptFeaturesxpsr Dedu.cornell.cs.nlp.spf.parser.ccg.features.basic.RuleUsageFeatureSet�k�d�L2� D scaleZ unaryRulesOnlyL 	ignoreSetq ~ xp?������� sr java.util.HashSet�D�����4  xpw   ?@      xsr Ledu.cornell.cs.nlp.spf.parser.ccg.features.basic.DynamicWordSkippingFeatures%�q�� L emptyCategoryq ~�L 
featureTagq ~ xpsq ~�p    sq ~$zT�lq ~&t EMPTYt DYNSKIPxq ~ sq ~ sq ~ 9   w   q ~ xq ~�sr %java.util.Collections$UnmodifiableSet��я��U  xq ~ sq ~�w   ?@     sr .edu.cornell.cs.nlp.spf.base.hashvector.KeyArgs���]e.ɘ I hashCodeL arg1q ~ L arg2q ~ L arg3q ~ L arg4q ~ L arg5q ~ xp2Iݬq ~ t 
TMPDEFAULTpppsq ~�wzq ~ t XEMEDEFAULTpppsq ~�'��q ~ t 
LEXDEFAULTpppxsr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoredLexicon�>�"z L lexemesq ~ (L lexemesByTypeq ~ (L 	templatesq ~ (xpsq ~ 2?@     0w   @   +q ~ �sq ~�w   ?@     q ~�q ~�q ~ �xq ~�sq ~�w   ?@     q ~xq ~�xq ~lsq ~�w   ?@     q ~�q ~ rq ~&q ~�q ~]q ~dq ~�q ~exq ~ �sq ~�w   ?@     q ~ �xq ~ �sq ~�w   ?@     q ~|q ~q ~ �xq ~
sq ~�w   ?@     q ~�q ~q ~�q ~�xq ~ osq ~�w   ?@     q ~Jq ~�q ~ Axq ~<sq ~�w   ?@     q ~6xq ~ �sq ~�w   ?@     q ~�q ~�q ~ �xq ~�sq ~�w   ?@     q ~�xq ~ =sq ~�w   ?@     q ~ +xq ~�sq ~�w   ?@     q ~�q ~�xq ~Vsq ~�w   ?@     q ~Hxq ~(sq ~�w   ?@     q ~q ~8q ~Zq ~�q ~�q ~@q ~Rq ~�xq ~ �sq ~�w   ?@     q ~ �xq ~usq ~�w   ?@     q ~mxq ~sq ~�w   ?@     q ~�q ~xq ~�sq ~�w   ?@     q ~�xq ~ �sq ~�w   ?@     q ~ �xq ~�sq ~�w   ?@     q ~�q ~�q ~.xq ~�sq ~�w   ?@     q ~�xq ~ sq ~�w   ?@     q ~ �xq ~ �sq ~�w   ?@     q ~ �xq ~sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~~sq ~�w   ?@     q ~vxq ~&sq ~�w   ?@     q ~xq ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~sq ~�w   ?@     q ~xq ~sq ~�w   ?@     q ~xq ~Zsq ~�w   ?@     q ~q ~Rxq ~�sq ~�w   ?@     q ~�xq ~zsq ~�w   ?@     q ~oq ~�q ~�xq ~msq ~�w   ?@     q ~0q ~�q ~�q ~(q ~bq ~nq ~�xq ~>sq ~�w   ?@     q ~�q ~�q ~3xq ~Esq ~�w   ?@     q ~?xq ~sq ~�w   ?@     q ~xq ~`sq ~�w   ?@     q ~Xxq ~1sq ~�w   ?@     q ~�q ~+q ~�q ~�xq ~ �sq ~�w   ?@     q ~ �q ~Hxq ~Gsq ~�w   ?@     q ~Axxsq ~ 2?@     w      q ~sq ~�w   ?@     q ~q ~�xq ~�sq ~�w   ?@     q ~�q ~|q ~�q ~Rq ~�q ~Jq ~�xq ~ �sq ~�w    ?@     q ~8q ~(q ~3q ~dq ~�q ~ �q ~q ~q ~�q ~eq ~Hq ~ �q ~�q ~ �q ~�q ~ �xq ~wsq ~�w   ?@     q ~�q ~oq ~�q ~�q ~ �xq ~�sq ~�w    ?@     q ~�q ~�q ~�q ~�q ~�q ~6q ~q ~�q ~q ~�q ~�q ~ +q ~?q ~+q ~q ~Aq ~ �q ~�q ~�xq ~%sq ~�w   ?@     q ~q ~bq ~�xq ~ �sq ~�w   ?@     q ~ �q ~ Axq ~ssq ~�w   ?@     q ~Zq ~]q ~nxq ~�sq ~�w   ?@     q ~�q ~�q ~q ~q ~vq ~�q ~�q ~mq ~xq ~�q ~Rq ~.xq ~�sq ~�w   ?@     q ~�q ~�q ~�q ~�q ~Xq ~�q ~Hq ~ �q ~�q ~�q ~ �xq ~�sq ~�w   ?@     q ~0q ~ rq ~�q ~�q ~�xq ~Esq ~�w   ?@     q ~�q ~&q ~@xxsq ~ 2?@     w      q ~�sq ~�w   ?@     q ~�q ~�xq ~�sq ~�w   ?@     q ~�q ~�q ~qxq ~�sq ~�w   ?@     q ~�q ~�q ~�q ~9xq ~ sq ~�w   ?@     q ~q ~*xq ~�sq ~�w   ?@     q ~�q ~iq ~`q ~�q ~�q ~�xq ~sq ~�w   ?@     q ~xq ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~%sq ~�w   ?@     q ~ xq ~{sq ~�w   ?@     q ~vq ~5xq ~Osq ~�w   ?@     q ~Jq ~�xq ~Vsq ~�w   ?@     q ~Qxxsr 9edu.cornell.cs.nlp.spf.base.hashvector.FastTreeHashVector;��tQ57� L valuest 0Lit/unimi/dsi/fastutil/objects/Object2DoubleMap;xpsr 5it.unimi.dsi.fastutil.objects.Object2DoubleAVLTreeMap�7y�J| I countL storedComparatort Ljava/util/Comparator;xr <it.unimi.dsi.fastutil.objects.AbstractObject2DoubleSortedMap�c����  xr 6it.unimi.dsi.fastutil.objects.AbstractObject2DoubleMap�o��K<z  xr ;it.unimi.dsi.fastutil.objects.AbstractObject2DoubleFunction�o��K<z D defRetValuexp          .psq ~�WD�t DYNSKIPppppw��      sq ~�W�"�q ~ t LEXt 0t 0pw        sq ~�W�#�q ~ q ~2t 0t 6pw@$      sq ~�W�&�q ~ q ~2t 1t 0pw@$      sq ~�W�&�q ~ q ~2t 1t 1pw����!asq ~�W�'Rq ~ q ~2t 1t 6pw��G:��f�sq ~�W�iq ~ q ~2t 10t 0pw        sq ~�W�iDq ~ q ~2t 10t 2pw@9�y��_sq ~�W�$�q ~ q ~2t 11t 11pw@7_��n�Ysq ~�W�%�q ~ q ~2t 11t 17pw        sq ~�W�(�q ~ q ~2t 11t 21pw@)�k��}sq ~�W�m�q ~ q ~2t 11t 8pw@3	�Wf�sq ~�W�,:q ~ q ~2t 12t 20pw@%��gi�fsq ~�W�qq ~ q ~2t 12t 4pw        sq ~�W�,xq ~ q ~2t 13t 12pw        sq ~�W�,�q ~ q ~2t 13t 16pw@5�~�B�sq ~�W�09q ~ q ~2t 14t 12pw@$      sq ~�W�0�q ~ q ~2t 14t 16pw?�Ԃ'6��sq ~�W�4q ~ q ~2t 15t 13pw@5oz�G�sq ~�W�48q ~ q ~2t 15t 14pw@5oz�G�sq ~�W�8q ~ q ~2t 16t 15pw@$      sq ~�W�;|q ~ q ~2t 17t 12pw@$      sq ~�W�;�q ~ q ~2t 17t 16pw?��ῶ��sq ~�Wć-q ~ q ~2t 18t 1pw@5oz�G�sq ~�Wć�q ~ q ~2t 18t 6pw        sq ~�Wċ�q ~ q ~2t 19t 6pw@4��`FX�sq ~�W�*xq ~ q ~2t 2t 1pw@6"S�.sq ~�W�*�q ~ q ~2t 2t 2pw        sq ~�WŖNq ~ q ~2t 20t 18pw        sq ~�WřUq ~ q ~2t 20t 22pw@$      sq ~�Wřtq ~ q ~2t 21t 13pw        sq ~�WŜ�q ~ q ~2t 21t 21pw@$      sq ~�WŜ�q ~ q ~2t 22t 10pw@$      sq ~�Wš�q ~ q ~2t 23t 19pw@5oz�G�sq ~�WŤZq ~ q ~2t 24t 10pw@$      sq ~�W��q ~ q ~2t 24t 5pw        sq ~�W��*q ~ q ~2t 25t 0pw@$      sq ~�W��Iq ~ q ~2t 25t 1pw��������sq ~�W��hq ~ q ~2t 25t 2pw���+�V�sq ~�W���q ~ q ~2t 25t 6pw��$J�F�sq ~�WŬ�q ~ q ~2t 26t 16pw@5�3̌�sq ~�Wų�q ~ q ~2t 27t 24pw@5�~�B�sq ~�W���q ~ q ~2t 27t 7pw        sq ~�W��q ~ q ~2t 28t 5pw@5�~�B�sq ~�W���q ~ q ~2t 29t 5pw?�Ԃ'5*�sq ~�W� Eq ~ q ~2t 29t 9pw@$      sq ~�W�.Xq ~ q ~2t 3t 2pw@1�g�s\�sq ~�W�.�q ~ q ~2t 3t 6pw��G>M�}�sq ~�W��q ~ q ~2t 30t 24pw@5�3̌�sq ~�W�R�q ~ q ~2t 30t 7pw        sq ~�W�U�q ~ q ~2t 31t 2pw@%���n�sq ~�W�V?q ~ q ~2t 31t 6pw        sq ~�W�Nq ~ q ~2t 32t 19pw@6z��sq ~�W�q ~ q ~2t 33t 23pw@$      sq ~�W�Tq ~ q ~2t 34t 15pw@$      sq ~�W� �q ~ q ~2t 35t 24pw?��ῶ��sq ~�W�ebq ~ q ~2t 35t 7pw@$      sq ~�W�!3q ~ q ~2t 36t 18pw@$      sq ~�W�$:q ~ q ~2t 36t 22pw        sq ~�W�(q ~ q ~2t 37t 23pw@$      sq ~�W�p)q ~ q ~2t 38t 3pw@$      sq ~�W�/�q ~ q ~2t 39t 25pw@$      sq ~�W�28q ~ q ~2t 4t 3pw@$      sq ~�WƁ�q ~ q ~2t 40t 20pw��ٴr	�sq ~�W�Ɵq ~ q ~2t 40t 4pw@5oz�G�sq ~�WƆ1q ~ q ~2t 41t 25pw@$      sq ~�Wƅ�q ~ q ~2t 42t 13pw@�߬~�lsq ~�WƆoq ~ q ~2t 42t 17pw        sq ~�WƊnq ~ q ~2t 43t 19pw?�v��+Sesq ~�WƐ�q ~ q ~2t 44t 20pw?]\��ʀ sq ~�W�գq ~ q ~2t 44t 4pw?�v��+Sesq ~�W���q ~ q ~2t 45t 0pw        sq ~�W��q ~ q ~2t 45t 1pw?�v��+Sesq ~�Wƕ�q ~ q ~2t 46t 19pw?�U(Osq ~�W���q ~ q ~2t 47t 1pw?�d��	sq ~�W��$q ~ q ~2t 47t 6pw        sq ~�WƟ�q ~ q ~2t 48t 20pw����o��sq ~�W��q ~ q ~2t 48t 4pw?��R��sq ~�WƟ�q ~ q ~2t 49t 11pw@�QC͊sq ~�WƠ:q ~ q ~2t 49t 13pw���}��sq ~�Wƣ�q ~ q ~2t 49t 21pw���'����sq ~�W���q ~ q ~2t 49t 8pw@��r�Q(sq ~�W�6q ~ q ~2t 5t 4pw@6u}Y��sq ~�W�:�q ~ q ~2t 50t 0pw        sq ~�W�:�q ~ q ~2t 50t 2pw�h:	
�msq ~�W�;<q ~ q ~2t 50t 6pw@���JJsq ~�W��Kq ~ q ~2t 51t 19pw?�L�O�Lsq ~�W���q ~ q ~2t 52t 20pw���v��sq ~�W�B�q ~ q ~2t 52t 4pw?��&�\�sq ~�W��q ~ q ~2t 53t 21pw?��v�Ecsq ~�W��q ~ q ~2t 54t 13pw?���B�Ssq ~�W�Wq ~ q ~2t 54t 21pw        sq ~�W��q ~ q ~2t 55t 13pw?���B�Ssq ~�W�	q ~ q ~2t 55t 21pw        sq ~�W�
q ~ q ~2t 56t 19pw        sq ~�W�q ~ q ~2t 57t 13pw?����l.�sq ~�W��q ~ q ~2t 57t 17pw        sq ~�W��q ~ q ~2t 58t 11pw?����c~ssq ~�W��q ~ q ~2t 58t 13pw?��}��=1sq ~�W�Y�q ~ q ~2t 58t 8pw?�[TM��ksq ~�W�Sq ~ q ~2t 59t 19pw?����sq ~�W�9�q ~ q ~2t 6t 5pw@5�3̌�sq ~�W�:tq ~ q ~2t 6t 9pw        sq ~�W�j�q ~ q ~2t 60t 21pw?��]=ްRsq ~�W�j�q ~ q ~2t 61t 13pw?��,7W�sq ~�WƳ�q ~ q ~2t 61t 8pw        sq ~�W�okq ~ q ~2t 62t 19pw?����Gsq ~�W�s,q ~ q ~2t 63t 19pw?��v���sq ~�Wƽ�q ~ q ~2t 64t 0pw��o��@h'sq ~�Wƾq ~ q ~2t 64t 1pw��t��vsq ~�Wƾ#q ~ q ~2t 64t 2pw?�E'�hsq ~�W�z�q ~ q ~2t 65t 19pw?��b�ȡQsq ~�Wǁ8q ~ q ~2t 66t 21pw?����v�sq ~�WǄ�q ~ q ~2t 67t 20pw@���ŏ�sq ~�W�ɤq ~ q ~2t 67t 4pw�����sq ~�Wǈ�q ~ q ~2t 68t 21pw        sq ~�W���q ~ q ~2t 68t 8pw@���ŏ�sq ~�Wǉ�q ~ q ~2t 69t 19pw?"��@ sq ~�W��Lq ~ q ~2t 7t 24pw?�Ԃ'6��sq ~�W�=�q ~ q ~2t 7t 7pw@$      sq ~�W���q ~ q ~2t 70t 20pw?����sq ~�W��q ~ q ~2t 71t 20pw?��)H��sq ~�W�'}q ~ q ~2t 71t 4pw        sq ~�W��tq ~ q ~2t 72t 20pw?��=��sq ~�W�+>q ~ q ~2t 72t 4pw        sq ~�W��q ~ q ~2t 73t 19pw?����Nsq ~�W�2�q ~ q ~2t 74t 2pw@����^sq ~�W�2�q ~ q ~2t 74t 6pw��^��Ov�sq ~�W��3q ~ q ~2t 75t 24pw        sq ~�W�6�q ~ q ~2t 75t 7pw?�99���sq ~�W��q ~ q ~2t 76t 25pw?�99���sq ~�W���q ~ q ~2t 77t 12pw?�99���sq ~�W�A�q ~ q ~2t 78t 3pw?�99���sq ~�W�E�q ~ q ~2t 79t 5pw        sq ~�W�F q ~ q ~2t 79t 9pw?�99���sq ~�W��-q ~ q ~2t 8t 13pw        sq ~�W���q ~ q ~2t 8t 17pw@$      sq ~�W�A�q ~ q ~2t 8t 8pw        sq ~�WǗ�q ~ q ~2t 80t 0pw?�$'��@sq ~�WǗ�q ~ q ~2t 80t 1pw��C��;�sq ~�WǗ�q ~ q ~2t 80t 2pw��:Uf��sq ~�W�S�q ~ q ~2t 81t 15pw?�99���sq ~�W�Woq ~ q ~2t 82t 13pw?�eo���sq ~�W�Z�q ~ q ~2t 82t 21pw�����97sq ~�WǠq ~ q ~2t 82t 8pw        sq ~�WǢ�q ~ q ~2t 83t 0pw        sq ~�Wǣq ~ q ~2t 83t 1pw���!�sq ~�Wǣ q ~ q ~2t 83t 2pw@�w�y#wsq ~�W�bUq ~ q ~2t 84t 20pw?�4[Y#losq ~�Wǧq ~ q ~2t 84t 4pw        sq ~�W�c.q ~ q ~2t 85t 17pw        sq ~�Wǫ\q ~ q ~2t 85t 8pw?��a� �sq ~�W�f5q ~ q ~2t 86t 11pw?�ȫ�
E�sq ~�W�f�q ~ q ~2t 86t 17pw        sq ~�W�j4q ~ q ~2t 87t 13pw?����/��sq ~�W�m�q ~ q ~2t 87t 21pw��[.�J,sq ~�Wǲ�q ~ q ~2t 87t 8pw        sq ~�W���q ~ q ~2t 9t 10pw        sq ~�W�E;q ~ q ~2t 9t 5pw?��ῶ��sq ~�W�E�q ~ q ~2t 9t 9pw@$      q ~�w?�      sq ~�e��q ~ t TMPt 0ppw?�VU���qsq ~�e���q ~ q ~	t 1ppw������y�sq ~�e�A>q ~ q ~	t 10ppw        sq ~�e�D�q ~ q ~	t 11ppw@��visq ~�e�H�q ~ q ~	t 12ppw?�()�sq ~�e�L�q ~ q ~	t 13ppw?���t�1Ysq ~�e�PBq ~ q ~	t 14ppw        sq ~�e�Tq ~ q ~	t 15ppw?�()�sq ~�e�W�q ~ q ~	t 16ppw?���
rFsq ~�e�[�q ~ q ~	t 17ppw        sq ~�e�_Fq ~ q ~	t 18ppw        sq ~�e�cq ~ q ~	t 19ppw?��N�3sq ~�e��q ~ q ~	t 2ppw@�s�V��sq ~�eص�q ~ q ~	t 20ppw?�3���]sq ~�eع^q ~ q ~	t 21ppw?�w͉d�sq ~�eؽq ~ q ~	t 22ppw        sq ~�e���q ~ q ~	t 23ppw        sq ~�e�ġq ~ q ~	t 24ppw?���
rFsq ~�e��bq ~ q ~	t 25ppw?�()�sq ~�e�Rq ~ q ~	t 3ppw?�()�sq ~�e�
q ~ q ~	t 4ppw?�0�l�Yssq ~�e��q ~ q ~	t 5ppw?���
rFsq ~�e��q ~ q ~	t 6ppw?�i_��sq ~�e�Vq ~ q ~	t 7ppw?�()�sq ~�e�q ~ q ~	t 8ppw@�� '�sq ~�e��q ~ q ~	t 9ppw?�()�q ~�w?�      sq ~�{H�q ~ t XEMEt 0ppw@$      sq ~�{H��q ~ q ~	Et 1ppw@#&|F�sq ~�{^�0q ~ q ~	Et 10ppw@9�y��_sq ~�{^��q ~ q ~	Et 11ppw@Aw-��]sq ~�{^��q ~ q ~	Et 12ppw@%��gi�fsq ~�{^�sq ~ q ~	Et 13ppw@$�y).sq ~�{^�4q ~ q ~	Et 14ppw@$Σ�v�sq ~�{_ �q ~ q ~	Et 15ppw@$      sq ~�{_�q ~ q ~	Et 16ppw@$      sq ~�{_wq ~ q ~	Et 17ppw@$��
���sq ~�{_8q ~ q ~	Et 18ppw@$      sq ~�{_�q ~ q ~	Et 19ppw@4��`FX�sq ~�{H��q ~ q ~	Et 2ppw@%SqKbsq ~�{_b�q ~ q ~	Et 20ppw@$      sq ~�{_fPq ~ q ~	Et 21ppw@$      sq ~�{_jq ~ q ~	Et 22ppw@$      sq ~�{_m�q ~ q ~	Et 23ppw@$      sq ~�{_q�q ~ q ~	Et 24ppw@$      sq ~�{_uTq ~ q ~	Et 25ppw@�Vޮ�Dsq ~�{_yq ~ q ~	Et 26ppw@$1qż�sq ~�{_|�q ~ q ~	Et 27ppw@$�y).sq ~�{_��q ~ q ~	Et 28ppw@$�y).sq ~�{_�Xq ~ q ~	Et 29ppw@$Σ�l�Jsq ~�{H�Dq ~ q ~	Et 3ppw@1���sq ~�{_��q ~ q ~	Et 30ppw@$1qż�sq ~�{_گq ~ q ~	Et 31ppw@%���n�sq ~�{_�pq ~ q ~	Et 32ppw@%U����	sq ~�{_�1q ~ q ~	Et 33ppw@$      sq ~�{_��q ~ q ~	Et 34ppw@$      sq ~�{_�q ~ q ~	Et 35ppw@$��
���sq ~�{_�tq ~ q ~	Et 36ppw@$      sq ~�{_�5q ~ q ~	Et 37ppw@$      sq ~�{_��q ~ q ~	Et 38ppw@$      sq ~�{_��q ~ q ~	Et 39ppw@$      sq ~�{H�q ~ q ~	Et 4ppw@$      sq ~�{`KMq ~ q ~	Et 40ppw@#12\oo�sq ~�{`Oq ~ q ~	Et 41ppw@$      sq ~�{`R�q ~ q ~	Et 42ppw@�߬~�lsq ~�{`V�q ~ q ~	Et 43ppw?�v��+Sesq ~�{`ZQq ~ q ~	Et 44ppw?֒�ǽ�Hsq ~�{`^q ~ q ~	Et 45ppw?�v��$9sq ~�{`a�q ~ q ~	Et 46ppw?�U(Osq ~�{`e�q ~ q ~	Et 47ppw?�d��	sq ~�{`iUq ~ q ~	Et 48ppw��i�Mǚsq ~�{`mq ~ q ~	Et 49ppw@+����Ssq ~�{H��q ~ q ~	Et 5ppw@%U�'V�"sq ~�{`��q ~ q ~	Et 50ppw@볬��sq ~�{`�mq ~ q ~	Et 51ppw?�L�O�Lsq ~�{`�.q ~ q ~	Et 52ppw?� �PvRsq ~�{`��q ~ q ~	Et 53ppw?��v�Ecsq ~�{`ΰq ~ q ~	Et 54ppw?���B�Ssq ~�{`�qq ~ q ~	Et 55ppw?���B�Ssq ~�{`�2q ~ q ~	Et 56ppw        sq ~�{`��q ~ q ~	Et 57ppw?����l.�sq ~�{`ݴq ~ q ~	Et 58ppw@ۤ˶Ksq ~�{`�uq ~ q ~	Et 59ppw?����sq ~�{H��q ~ q ~	Et 6ppw@$1qż�sq ~�{a4q ~ q ~	Et 60ppw?��]=�¤sq ~�{a7�q ~ q ~	Et 61ppw?��,7W�sq ~�{a;�q ~ q ~	Et 62ppw?����Gsq ~�{a?Nq ~ q ~	Et 63ppw?��v���sq ~�{aCq ~ q ~	Et 64ppw���\'���sq ~�{aF�q ~ q ~	Et 65ppw?��b�ȡQsq ~�{aJ�q ~ q ~	Et 66ppw?����v�sq ~�{aNRq ~ q ~	Et 67ppw?����v�sq ~�{aRq ~ q ~	Et 68ppw@���4QNsq ~�{aU�q ~ q ~	Et 69ppw?"��@ sq ~�{H�Hq ~ q ~	Et 7ppw@$Σ�v�sq ~�{a�jq ~ q ~	Et 70ppw?����sq ~�{a�+q ~ q ~	Et 71ppw?��)H��sq ~�{a��q ~ q ~	Et 72ppw?��=��sq ~�{a��q ~ q ~	Et 73ppw?����Nsq ~�{a�nq ~ q ~	Et 74ppw@;��Esq ~�{a�/q ~ q ~	Et 75ppw?�99���sq ~�{a��q ~ q ~	Et 76ppw?�99���sq ~�{a±q ~ q ~	Et 77ppw?�99���sq ~�{a�rq ~ q ~	Et 78ppw?�99���sq ~�{a�3q ~ q ~	Et 79ppw?�99���sq ~�{H�	q ~ q ~	Et 8ppw@$      sq ~�{b�q ~ q ~	Et 80ppw��>��W��sq ~�{b �q ~ q ~	Et 81ppw?�99���sq ~�{b$Kq ~ q ~	Et 82ppw?�ȫ�
F�sq ~�{b(q ~ q ~	Et 83ppw?��a�!Qsq ~�{b+�q ~ q ~	Et 84ppw?�4[Y#?sq ~�{b/�q ~ q ~	Et 85ppw?��a� �sq ~�{b3Oq ~ q ~	Et 86ppw?�ȫ�
E�sq ~�{b7q ~ q ~	Et 87ppw?��a��sq ~�{H��q ~ q ~	Et 9ppw@$��
�{Sq ~�w?�      sq ~���#)t LOGEXPt CPP1q ~q ~ �q ~ �w��G>M�}�sq ~�1��q ~	�q ~	�q ~q ~�q ~ �w��FJ�I/+sq ~�d��q ~	�q ~	�q ~q ~ �q ~ �w��A#��Asq ~�6X�{q ~	�q ~	�q ~q ~ �q ~ �w?�C����sq ~��Z��q ~	�q ~	�q ~q ~ �q ~�w?��k�j�*sq ~�V�b�q ~	�q ~	�q ~q ~Oq ~ �w��,L�#Basq ~�(��-q ~	�q ~	�q ~q ~Oq ~ �w@���Y��sq ~���`�q ~	�q ~	�q ~q ~Oq ~�w?�f�v��sq ~��=�,q ~	�q ~	�q ~q ~Oq ~ �w���JM�hmsq ~�gGE�q ~	�q ~	�q ~q ~Oq ~�w?����sq ~���l�q ~	�q ~	�q ~q ~q ~w?��
�i�sq ~�Q���q ~	�q ~	�q ~q ~q ~ �w@YA���sq ~׾�&�q ~	�q ~	�q ~q ~q ~ �w?�BX�/\+sq ~�I�vDq ~	�q ~	�q ~q ~q ~�w?����sq ~�D��q ~	�q ~	�q ~q ~q ~Ow@�k�을sq ~�G٢0q ~	�t REPTq ~q ~ �pw����|��sq ~��<agq ~	�q ~
q ~q ~�pw��@'͵�sq ~�r��q ~	�q ~
q ~q ~ �pw���;�.7�sq ~�d!+�t RULEt <applypppw?�A�fSPsq ~׌�	�q ~
t >applypppw@%Pd=lG�sq ~�"A�q ~
t >comp1pppw��9~�J<sq ~�4::�q ~
t 	>thatlesspppw��l���fsq ~�Z�q ~
t >trcomp1pppw?���Y8ىsq ~�Կq ~
t lexpppw@)���Ӄsq ~�R롞q ~
t shift_pppppw?�O�dm-*x