�� sr -edu.cornell.cs.nlp.spf.parser.ccg.model.Model�5B��B�~ L featureSetst Ljava/util/List;L independentLexicalFeatureSetsq ~ L invalidFeaturest Ljava/util/Set;L lexicont -Ledu/cornell/cs/nlp/spf/ccg/lexicon/ILexicon;L thetat 4Ledu/cornell/cs/nlp/spf/base/hashvector/IHashVector;xpsr &java.util.Collections$UnmodifiableList�%1�� L listq ~ xr ,java.util.Collections$UnmodifiableCollectionB ��^� L ct Ljava/util/Collection;xpsr java.util.LinkedList)S]J`�"  xpw   sr Pedu.cornell.cs.nlp.spf.parser.ccg.factoredlex.features.FactoredLexicalFeatureSet�g�պ��� D 
entryScaleI lexemeNextIdD lexemeScaleI nonFactoredNextIdI templateNextIdD templateScaleL entryInitialScorert :Ledu/cornell/cs/nlp/utils/collections/ISerializableScorer;L 	lexemeIdst 5Lit/unimi/dsi/fastutil/objects/Object2IntOpenHashMap;L lexemeInitialScorerq ~ L nonFactoredIdsq ~ L templateIdsq ~ L templateInitialScorerq ~ xr Iedu.cornell.cs.nlp.spf.parser.ccg.model.lexical.AbstractLexicalFeatureSetZ���n3�� Z computeSyntaxAttributeFeaturesL 
featureTagt Ljava/lang/String;L ignoreFiltert Ljava/util/function/Predicate;xp t FACLEXsr !java.lang.invoke.SerializedLambdaoaД,)6� 
I implMethodKind[ capturedArgst [Ljava/lang/Object;L capturingClasst Ljava/lang/Class;L functionalInterfaceClassq ~ L functionalInterfaceMethodNameq ~ L "functionalInterfaceMethodSignatureq ~ L 	implClassq ~ L implMethodNameq ~ L implMethodSignatureq ~ L instantiatedMethodTypeq ~ xp   ur [Ljava.lang.Object;��X�s)l  xp    vr 0edu.cornell.cs.nlp.utils.function.PredicateUtils           xpt java/util/function/Predicatet testt (Ljava/lang/Object;)Zt 0edu/cornell/cs/nlp/utils/function/PredicateUtilst lambda$alwaysTrue$bcad8f2c$1q ~ q ~ ?�         n?�             ?�������sr Eedu.cornell.cs.nlp.spf.parser.ccg.features.basic.scorer.UniformScorerQ�B���S D scorexp        sr 3it.unimi.dsi.fastutil.objects.Object2IntOpenHashMap         F fI sizexr 3it.unimi.dsi.fastutil.objects.AbstractObject2IntMap�o��K<z  xr 8it.unimi.dsi.fastutil.objects.AbstractObject2IntFunction�o��K<z I defRetValuexp    ?@     nsr 9edu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.Lexeme	I����� I hashCodeCacheL 
attributesq ~ L 	constantsq ~ L 
propertiest Ljava/util/Map;L 	signaturet GLedu/cornell/cs/nlp/spf/ccg/lexicon/factored/lambda/FactoringSignature;L tokenst ,Ledu/cornell/cs/nlp/spf/base/token/TokenSeq;xp��g�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sr 0edu.cornell.cs.nlp.spf.mr.lambda.LogicalConstant=Q��� L baseNameq ~ L nameq ~ xr %edu.cornell.cs.nlp.spf.mr.lambda.Term�(G^� L typet .Ledu/cornell/cs/nlp/spf/mr/language/type/Type;xr 2edu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression
n�tL�h  xpsr 3edu.cornell.cs.nlp.spf.mr.language.type.ComplexType� �g��V L domainq ~ 2L rangeq ~ 2xr ,edu.cornell.cs.nlp.spf.mr.language.type.Typeg���� I hashCodeCacheL nameq ~ xp?z�t 	<e,<e,t>>sr 0edu.cornell.cs.nlp.spf.mr.language.type.TermType��6��ǭ L parentt 2Ledu/cornell/cs/nlp/spf/mr/language/type/TermType;xq ~ 6   et epsq ~ 5|-t <e,t>q ~ ;sq ~ 9   tt tpt neart near:<e,<e,t>>sq ~ 0q ~ =t agentt agent:<e,t>xq ~ /q ~ .sr %java.util.Collections$UnmodifiableMap��t�B L mq ~ (xpsq ~ Fsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t origint fixed_domainxsr Eedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoringSignature�ڝ�U鞉 I hashCodeI numAttributesL typesq ~ xp�W;    sq ~ sr java.util.ArrayListx����a� I sizexp   w   q ~ 7q ~ =xq ~ Qsr *edu.cornell.cs.nlp.spf.base.token.TokenSeq�py��An I hashCode[ tokenst [Ljava/lang/String;xp4P�ur [Ljava.lang.String;��V��{G  xp   t movet tow   sq ~ '��3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~ ]q ~ \sq ~ Fsq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kt genlexxsq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~ esq ~ R 3�1uq ~ U   t nextw   5sq ~ '~�_q ~ ,sq ~ sq ~ sq ~ 
w   q ~ Cxq ~ lq ~ ksq ~ Fq ~ Hsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~ pq ~ Tw   sq ~ '��
sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 7t rightt right:<e,<e,t>>q ~ Cxq ~ uq ~ tsq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~ }sq ~ R��uq ~ U   t standw   6sq ~ '{�%sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ vq ~ Cxq ~ �q ~ �sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~ �sq ~ R $�/uq ~ U   t Movew   9sq ~ '�m�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ vq ~ Cxq ~ �q ~ �sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~ �sq ~ Rzj�uq ~ U   t robotw   Esq ~ 'H׫sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ =t blockt block:<e,t>xq ~ �q ~ �sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~ �sq ~ R 3�1uq ~ U   q ~ hw   >sq ~ '�b�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~ �q ~ �sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~ �sq ~ R���uq ~ U   q ~ �w   sq ~ ' 8)Csq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~ �sq ~ R 7�uq ~ U   t withw   dsq ~ ' 4psq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~ �sq ~ R 3�1uq ~ U   q ~ hw   Tsq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~ �sq ~ R  �uq ~ U   q ~ Xw    sq ~ '�@�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M  �    sq ~ sq ~ P    w    xq ~ �sq ~ R�@(uq ~ U   t pleasew   sq ~ 'A+�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 7t leftt left:<e,<e,t>>xq ~ �q ~ �sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~ �sq ~ R 2�Euq ~ U   q ~ �w   sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~sq ~ R  cuq ~ U   t inw   Qsq ~ ' +�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~
sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M  �    sq ~ sq ~ P    w    xq ~sq ~ R �Muq ~ U   t putw   sq ~ '��x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~sq ~ R�� Huq ~ U   t Pleasew   ?sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~&q ~%sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~+sq ~ R  �uq ~ U   t byw   Osq ~ '�%�Ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~3q ~2sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~9sq ~ Rg�Wuq ~ U   q ~ Wq ~ Aw   sq ~ '־-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~@q ~?sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~Esq ~ R �uq ~ U   t Enterw   msq ~ '  �(sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~Mq ~Lsq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~Rsq ~ R  �uq ~ U   t Dow   <sq ~ 'C%�q ~0sq ~ sq ~ sq ~ 
w   q ~ 4xq ~Yq ~Xsq ~ Fq ~5sq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~]q ~:w   sq ~ 'z��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~bq ~asq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~gsq ~ Rzj�uq ~ U   q ~ �w   Jsq ~ 'X��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ =t redt 	red:<e,t>xq ~nq ~msq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~vsq ~ R  �uq ~ U   t mew   bsq ~ 'Ҿ%�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~~q ~}sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R  �uq ~ U   q ~ Xw   &sq ~ 's���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ =t roomt 
room:<e,t>xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R8��uq ~ U   t coloredw   ,sq ~ '<�Ըsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~�sq ~ R 3�fuq ~ U   q ~ Aw   sq ~ '͖Y)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 7q ~t in:<e,<e,t>>q ~ Cxq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R4P�uq ~ U   q ~ Wq ~ Xw   sq ~ '�FĘsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~�sq ~ R  cuq ~ U   q ~w   sq ~ '�)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R �Uuq ~ U   t farw   Zsq ~ 'w�(sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Cxq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R �suq ~ U   t goq ~ Xw   sq ~ ' 0�nsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R 0R/uq ~ U   t cant youw   	sq ~ ' �Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R zuq ~ U   t andw   ^sq ~ 'ׅ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R���uq ~ U   t Standw   \sq ~ ' 3�Nsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~sq ~ R 3<uq ~ U   q ~ Ww   /sq ~ '�<Ssq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~sq ~ R��uq ~ U   q ~ �w   $sq ~ 'B�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~q ~sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~%sq ~ R=��uq ~ U   q ~ hq ~ Xw   sq ~ '_D�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~,q ~+sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~1sq ~ Rw�Zuq ~ U   q ~ ww   7sq ~ '�HY�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~8q ~7sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~>sq ~ R �suq ~ U   q ~�q ~ Xw   sq ~ 'rK�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ =t doort 
door:<e,t>xq ~Eq ~Dsq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~Nsq ~ R /#�uq ~ U   q ~Gw   sq ~ ' 6qsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~Uq ~Tsq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~Zsq ~ R 5�@uq ~ U   t spotw   Gsq ~ '�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~bq ~asq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~hsq ~ R 1f�uq ~ U   t intow   
sq ~ '�߁sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~pq ~osq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~usq ~ R !juq ~ U   t Findw   lsq ~ ' �sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~}q ~|sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R �Uuq ~ U   q ~�w   isq ~ '+�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R0l��uq ~ U   t Positionw   esq ~ 'Y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R 7�uq ~ U   q ~ �w   gsq ~ ';_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R  �uq ~ U   q ~ Xw   0sq ~ '�w�Ysq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R�w�uq ~ U   t towardsw   `sq ~ '��Ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R 3<uq ~ U   q ~ Ww   Usq ~ '�B{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R 5ݕuq ~ U   t sidew   Rsq ~ '�Vusq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R��6uq ~ U   t closew   Wsq ~ '��Bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R  uq ~ U   t ofw   4sq ~ ';��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R 5�uq ~ U   q ~�w   sq ~ 'X�h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~ q ~�w   Vsq ~ '�?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ vq ~ Cxq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~
sq ~ R 3<uq ~ U   q ~ Ww   Csq ~ '  x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~sq ~ R   �uq ~ U   t aw   Fsq ~ '��s'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ Cxq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~#sq ~ Rzj�uq ~ U   q ~ �w   *sq ~ '  �\sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~*q ~)sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~/sq ~ R  uq ~ U   t onw   ]sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~7q ~6sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~<sq ~ R  �uq ~ U   t sow   Ksq ~ '�{�q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~Cq ~Bsq ~ Fq ~�sq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~Gq ~�w   sq ~ '�u0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~Lq ~Ksq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~Qsq ~ R��uq ~ U   t chairw   "sq ~ '�c��q ~5sq ~ sq ~ sq ~ 
w   q ~�q ~ Cxq ~Xq ~Wsq ~ Fq ~:sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~\q ~?w   sq ~ ''�Ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ Cxq ~aq ~`sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~fsq ~ RPŴ�uq ~ U   t Proceedw   ;sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~nq ~msq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~ssq ~ R  huq ~ U   t isw   Msq ~ ' 3?sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~{q ~zsq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R 2��uq ~ U   t lookw   _sq ~ '<�X�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~�sq ~ R  �uq ~ U   q ~.w   sq ~ 'B��q ~ ,sq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Fq ~ Hsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~�q ~ Tw   sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ vq ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R���uq ~ U   q ~w   Asq ~ 'ǕD�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R 3<uq ~ U   q ~ Ww   @sq ~ 'V�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R�� Huq ~ U   q ~!w   .sq ~ '}g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Cxq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R�CCuq ~ U   q ~ Dw    sq ~ '�BFsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R 5�uq ~ U   q ~�w   Isq ~ 'X��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�q ~�w   3sq ~ 'Y�>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R 5ݕuq ~ U   q ~�w   Xsq ~ '^p��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R��uq ~ U   q ~Tw   Ysq ~ '���1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~sq ~ R $�/uq ~ U   q ~ �w   %sq ~ 'ǆ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ Cxq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~q ~w   'sq ~ '0mu�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~sq ~ R0l��uq ~ U   q ~�w   Dsq ~ '  �zsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~#sq ~ R  ;uq ~ U   t hew   Lsq ~ '�e�)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~+q ~*sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~0q ~�w   +sq ~ ' 8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~5q ~4sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M  �    sq ~ sq ~ P    w    xq ~;sq ~ R ��uq ~ U   t thew   sq ~ 'f��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ vq ~ Cxq ~Cq ~Bsq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~Hsq ~ RRP��uq ~ U   t 
positionedw   Nsq ~ 'l�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ =t greent green:<e,t>xq ~Pq ~Osq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~Ysq ~ R��Auq ~ U   q ~Rw   sq ~ '  �Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~`q ~_sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~esq ~ R  uq ~ U   q ~�w   !sq ~ '~H3q ~0sq ~ sq ~ sq ~ 
w   q ~ Cxq ~kq ~jsq ~ Fq ~5sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~oq ~:w   sq ~ '�b8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ Cxq ~tq ~ssq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~yq ~�w   (sq ~ 'J��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ =t bluet 
blue:<e,t>xq ~~q ~}sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R .0�uq ~ U   q ~�w   sq ~ '%�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�q ~Iw   [sq ~ 'Ҿ Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R  	Fuq ~ U   t Gow   Psq ~ ' %(nsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R $�/uq ~ U   q ~ �w   sq ~ ' 6U�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R 5ݕuq ~ U   q ~�w   2sq ~ 'x:�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ Rw�Zuq ~ U   q ~ ww   fsq ~ '�L3sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R���uq ~ U   q ~w   1sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R  	Fuq ~ U   q ~�w   #sq ~ 'XΖxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~ R ��uq ~ U   q ~pw   sq ~ 'ҿ�uq ~�sq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~�q ~�sq ~ Fq ~�sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�q ~�w   sq ~ ' 1��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~ R 1f�uq ~ U   q ~kw   Bsq ~ ' 5�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~sq ~ R 5�uq ~ U   q ~�w   csq ~ 'Y_]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~oxq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~sq ~ R 4��uq ~ U   t pinkw   -sq ~ ' #Psq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fsq ~ Fq ~ `sq ~ M  �    sq ~ sq ~ P    w    xq ~ sq ~ R �uq ~ U   t notw   =sq ~ '�DO1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~(q ~'sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~-sq ~ R 7�uq ~ U   q ~ �w   ksq ~ 'ҿ�Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~4q ~3sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~9q ~�w   jsq ~ '�`�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~>q ~=sq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~Cq ~2w   :sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~Hq ~Gsq ~ Fsq ~ Fq ~ `sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~Mq ~ww   asq ~ '�c�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~Rq ~Qsq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~Wsq ~ R��6uq ~ U   q ~�w   8sq ~ '�8��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~^q ~]sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~csq ~ Rzj�uq ~ U   q ~ �w   hsq ~ '�H�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~jq ~isq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~oq ~ ~w   Ssq ~ '�b�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ Cxq ~tq ~ssq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~yq ~�w   )sq ~ 'M��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ vxq ~~q ~}sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~�sq ~ Rw�Zuq ~ U   q ~ ww   sq ~ '<���q ~�sq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Fq ~�sq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~�q ~�w   sq ~ '�u��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ Cxq ~�q ~�sq ~ Fsq ~ Fq ~ `sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sq ~ R�z�uq ~ U   t Robotw   Hxsq ~ !        sq ~ #    ?@      xsq ~ #    ?@     sr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.LexicalTemplateg��%��	 I hashCodeL 	argumentsq ~ L 
propertiesq ~ (L 	signatureq ~ )L templatet 0Ledu/cornell/cs/nlp/spf/ccg/categories/Category;xp�*z5sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 7t #0<e,<e,t>>t #0<e,<e,t>>:<e,<e,t>>sq ~ 0q ~ =t #0<e,t>t #0<e,t>:<e,t>xq ~�q ~�sq ~ Fq ~5sq ~ M�W;    sq ~ sq ~ P   w   q ~ 7q ~ =xq ~�sr 5edu.cornell.cs.nlp.spf.ccg.categories.ComplexCategory�f�Ք�nl I hashCodeCacheL syntaxt <Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/ComplexSyntax;xr .edu.cornell.cs.nlp.spf.ccg.categories.CategorycK=�.A� L 	semanticst Ljava/lang/Object;xpsr 'edu.cornell.cs.nlp.spf.mr.lambda.Lambda��Kβ�� L argumentt +Ledu/cornell/cs/nlp/spf/mr/lambda/Variable;L bodyt 4Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L typet 5Ledu/cornell/cs/nlp/spf/mr/language/type/ComplexType;xq ~ 3sr )edu.cornell.cs.nlp.spf.mr.lambda.Variable�u#$rP L 	singletonq ~ xq ~ 1q ~ ;sr 5it.unimi.dsi.fastutil.objects.ReferenceSets$Singleton�7y�J| L elementq ~�xpq ~�sr (edu.cornell.cs.nlp.spf.mr.lambda.Literalŕtb��� [ 	argumentst 5[Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L 	predicateq ~�[ 	signaturet /[Ledu/cornell/cs/nlp/spf/mr/language/type/Type;L typeq ~ 2xq ~ 3ur 5[Ledu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression;|�㰢�[i  xp   sq ~�uq ~�   sq ~�sq ~�q ~ ;sq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�ur /[Ledu.cornell.cs.nlp.spf.mr.language.type.Type;>L5��  xp   q ~ ;q ~ ?sr 4it.unimi.dsi.fastutil.objects.ReferenceSets$EmptySet�7y�J|  xpq ~ =q ~�sq ~ 0sq ~ 5I:��t 	<<e,t>,e>q ~ =q ~ ;q ~>t the:<<e,t>,e>uq ~�   q ~ =q ~ ;q ~�q ~�q ~�uq ~�   q ~ ;q ~ ;q ~ ?q ~�q ~ =���.sr :edu.cornell.cs.nlp.spf.ccg.categories.syntax.ComplexSyntax$���q\P^ I hashCodeI 	numSlahesL leftt 5Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax;L rightq ~�L slasht 4Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Slash;xr 3edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntaxʊ�	�|��  xpȠU�   sr @edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntax$SimpleSyntax��eBg� I hashCodeL 	attributeq ~ L labelq ~ xq ~� 3�t nonet Ssq ~� 4�wq ~�t NPsr 2edu.cornell.cs.nlp.spf.ccg.categories.syntax.Slashѕ�����> C cxp /w   sq ~�(�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~�sq ~�sq ~�q ~ =sq ~�q ~�sq ~�sq ~�q ~ ;sq ~�q ~�sq ~�uq ~�   q ~�sr ;it.unimi.dsi.fastutil.objects.ReferenceSets$UnmodifiableSet�7y�J|  xr Iit.unimi.dsi.fastutil.objects.ReferenceCollections$UnmodifiableCollection�7y�J| L 
collectiont 3Lit/unimi/dsi/fastutil/objects/ReferenceCollection;xpsr 2it.unimi.dsi.fastutil.objects.ReferenceOpenHashSet         F fI sizexp?@     q ~�q ~�xq ~�uq ~�   q ~ ;q ~ ?sq ~�sq ~�?@     q ~�xq ~ =q ~�sq ~ 5JW`Lt <<e,t>,<e,t>>q ~ =q ~ =(�>sq ~��|��   q ~�q ~�q ~�w   sq ~��7�'sq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Fq ~�sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~sq ~�sq ~�sq ~�q ~ ;sq ~�q ~
sq ~�uq ~�   sq ~�uq ~�   sq ~�sq ~�q ~ ;sq ~�q ~sq ~�uq ~�   q ~q ~q ~�uq ~�   q ~ ;q ~ ?q ~�q ~ =q ~�q ~�uq ~�   q ~ =q ~ ;q ~
q ~q ~�uq ~�   q ~ ;q ~ ;q ~ ?q ~�q ~ =�).sq ~�ȠU�   q ~�q ~�q ~�w   
sq ~�(W~sq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Fq ~7sq ~ M  �    sq ~ sq ~ P    w    xq ~ sq ~�sq ~�sq ~�q ~ =sq ~�q ~#sq ~�sq ~�q ~ ;sq ~�q ~&sq ~�uq ~�   q ~&sq ~�sq ~�?@     q ~#q ~&xq ~#uq ~�   q ~ ;q ~ ?sq ~�sq ~�?@     q ~#xq ~ =q ~�q ~�(S�sq ~��z�M   sq ~� 3�kq ~�t Nq ~0q ~�w   sq ~��?kisq ~ sq ~ sq ~ 
w    xq ~5q ~4sq ~ Fq ~sq ~ M  �    sq ~ sq ~ P    w    xq ~9sq ~�sq ~�sq ~�q ~ ;sq ~�q ~<sq ~�sq ~�q ~ =sq ~�q ~?sq ~�uq ~�   q ~<sq ~�sq ~�?@     q ~<q ~?xq ~?uq ~�   q ~ ;q ~ ?sq ~�sq ~�?@     q ~<xsq ~ 5I:�et 	<<e,t>,t>q ~ =q ~ ?q ~�sq ~ 5e5}\t <e,<<e,t>,t>>q ~ ;q ~H�?g�sq ~�+���   sq ~�ȡ>Z   q ~�sq ~� 4��q ~�t PPq ~�q ~�q ~�w   	sq ~�t�,sq ~ sq ~ sq ~ 
w   q ~�xq ~Sq ~Rsq ~ Fq ~:sq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~Wsq ~�sq ~�sq ~�q ~ ;sq ~�q ~Zsq ~�uq ~�   sq ~�uq ~�   sq ~�sq ~�q ~ ;sq ~�q ~asq ~�uq ~�   q ~aq ~bq ~ Cuq ~�   q ~ ;q ~ ?q ~�q ~ =q ~�q ~�uq ~�   q ~ =q ~ ;q ~Zq ~[q ~�uq ~�   q ~ ;q ~ ;q ~ ?q ~�q ~ =t��sq ~�ȠU�   q ~�q ~�q ~�w   sq ~����sq ~ sq ~ sq ~ 
w    xq ~lq ~ksq ~ Fq ~ �sq ~ M  �    sq ~ sq ~ P    w    xq ~psq ~�sq ~�sq ~�q ~ ?sq ~�q ~sq ~sq ~�sq ~ 5��t <t,t>q ~ ?q ~ ?���sq ~��|�   q ~�q ~�sq ~� \w   sq ~�IH�xsq ~ sq ~ sq ~ 
w   q ~�xq ~|q ~{sq ~ Fq ~Usq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~�sq ~�sq ~�q ~ =sq ~�q ~�sq ~�sq ~�q ~ ;sq ~�q ~�sq ~�uq ~�   sq ~�uq ~�   q ~�q ~�q ~�uq ~�   q ~ ;q ~ ?sq ~�uq ~�   q ~�sq ~�sq ~�?@     q ~�q ~�xq ~�uq ~�   q ~ ;q ~ ?sq ~�sq ~�?@     q ~�q ~�xsq ~ 0sr <edu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType&��M
� I minArgsZ orderSensitiveL optiont ELedu/cornell/cs/nlp/spf/mr/language/type/RecursiveComplexType$Option;xq ~ 5l�6�t <t*,t>q ~ ?q ~ ?    sr Cedu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType$Option�^g� �� Z isOrderSensitiveI 
minNumArgsxp    q ~�t 
and:<t*,t>uq ~�   q ~ ?q ~ ?q ~ ?sq ~�sq ~�?@     q ~�xq ~ =q ~�q ~�R:L]sq ~��z�M   q ~0q ~0q ~�w    sq ~���'sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Fq ~ �sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sr 4edu.cornell.cs.nlp.spf.ccg.categories.SimpleCategory��4_C� I hashCodeCacheL syntaxt BLedu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax$SimpleSyntax;xq ~�sq ~�sq ~�q ~ ;sq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�uq ~�   q ~ ;q ~ ?q ~�q ~ =�Ǵq ~0w   sq ~�x�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fsq ~ Fsq ~ I?@     w      q ~ Kq ~ Lxsq ~ M  �    sq ~ sq ~ P    w    xq ~�sq ~�sq ~�sq ~�q ~ =sq ~�q ~�sq ~�uq ~�   sq ~�sq ~�q ~ ;sq ~�q ~�sq ~�uq ~�   q ~�sq ~�sq ~�?@     q ~�q ~�xq ~�uq ~�   q ~ ;q ~ ?sq ~�sq ~�?@     q ~�xq ~ =q ~�q ~�uq ~�   q ~ =q ~ ;q ~�q ~�x~'sq ~��ƥY   q ~�q ~0q ~�w   sq ~�'���sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Fq ~!sq ~ M?z��    sq ~ sq ~ P   w   q ~ 7xq ~�sq ~�sq ~�sq ~�q ~ ;sq ~�q ~�sq ~�sq ~�q ~ ;sq ~�q ~�sq ~�uq ~�   q ~�q ~�sq ~�sq ~�?@     q ~�q ~�xq ~�uq ~�   q ~ ;q ~ ;q ~ ?sq ~�sq ~�?@     q ~�xq ~ =q ~�q ~ 7':sq ~ԫR   sq ~��P�   q ~Nq ~�q ~�q ~�q ~xw   sq ~�󓠪sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Fq ~5sq ~ M|#    sq ~ sq ~ P   w   q ~ =xq ~�sq ~�sq ~�q ~�sq ~�uq ~�   sq ~�uq ~�   sq ~�q ~�sq ~�uq ~�   q ~�q ~�q ~�uq ~�   q ~ ;q ~ ?q ~�q ~ =q ~�q ~�uq ~�   q ~ =q ~ ;q ~�q ~�q ~ 4uq ~�   q ~ ;q ~ ;q ~ ?q ~�q ~ =��<�q ~�w   sq ~����sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Fq ~�sq ~ M  �    sq ~ sq ~ P    w    xq ~ sq ~�sq ~�sq ~�q ~ ?sq ~�q ~q ~q ~�q ~u���sq ~��|��   q ~�q ~�q ~�w   xsq ~ !        sr Yedu.cornell.cs.nlp.spf.parser.ccg.features.lambda.LogicalExpressionCoordinationFeatureSet�4tHWcg+ Z cpapFeaturesZ cpp1FeaturesZ reptFeaturesxpsr Dedu.cornell.cs.nlp.spf.parser.ccg.features.basic.RuleUsageFeatureSet�k�d�L2� D scaleZ unaryRulesOnlyL 	ignoreSetq ~ xp?�       sr java.util.HashSet�D�����4  xpw   ?@      xsr Ledu.cornell.cs.nlp.spf.parser.ccg.features.basic.DynamicWordSkippingFeatures%�q�� L emptyCategoryq ~�L 
featureTagq ~ xpsq ~�p    sq ~�zT�lq ~�t EMPTYt DYNSKIPsr Yedu.cornell.cs.nlp.spf.parser.ccg.features.lambda.LogicalExpressionCooccurrenceFeatureSetf��C �c�  xpxq ~ sq ~ sq ~ P   w   q ~ xq ~sr %java.util.Collections$UnmodifiableSet��я��U  xq ~ sq ~w   ?@     sr .edu.cornell.cs.nlp.spf.base.hashvector.KeyArgs���]e.ɘ I hashCodeL arg1q ~ L arg2q ~ L arg3q ~ L arg4q ~ L arg5q ~ xp2Iݬq ~ t 
TMPDEFAULTpppsq ~wzq ~ t XEMEDEFAULTpppsq ~'��q ~ t 
LEXDEFAULTpppxsr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoredLexicon�>�"z L lexemesq ~ (L lexemesByTypeq ~ (L 	templatesq ~ (xpsq ~ I?@     `w   �   8q ~sq ~w   ?@     q ~
xq ~ fsq ~w   ?@     q ~ Yq ~ �q ~ �xq ~gsq ~w   ?@     q ~]xq ~�sq ~w   ?@     q ~�q ~q ~�q ~ �xq ~!sq ~w   ?@     q ~xq ~Xsq ~w   ?@     q ~�q ~Nxq ~�sq ~w   ?@     q ~�xq ~fsq ~w   ?@     q ~�q ~\q ~�xq ~�sq ~w   ?@     q ~"q ~�xq ~Isq ~w   ?@     q ~?q ~�xq ~�sq ~w   ?@     q ~�q ~'xq ~=sq ~w   ?@     q ~3xq ~0sq ~w   ?@     q ~&xq ~sq ~w   ?@     q ~q ~ qq ~fxq ~�sq ~w   ?@     q ~@q ~ iq ~�q ~ +q ~�xq ~sq ~w   ?@     q ~xq ~�sq ~w   ?@     q ~�xq ~�sq ~w   ?@     q ~�q ~�q ~�xq ~Rsq ~w   ?@     q ~Hq ~�xq ~Zsq ~w   ?@     q ~Lxq ~�sq ~w   ?@     q ~�q ~�q ~�xq ~�sq ~w   ?@     q ~�q ~:q ~(q ~zxq ~<sq ~w   ?@     q ~1xq ~isq ~w   ?@     q ~^q ~�xq ~:sq ~w   ?@     q ~hq ~/q ~Vxq ~ �sq ~w   ?@     q ~$q ~�q ~ �xq ~�sq ~w   ?@     q ~�q ~�q ~�xq ~vsq ~w   ?@     q ~lxq ~�sq ~w   ?@     q ~zxq ~ �sq ~w   ?@     q ~zq ~�q ~ �q ~pxq ~$sq ~w   ?@     q ~xq ~sq ~w   ?@     q ~�q ~�q ~q ~xq ~�sq ~w   ?@     q ~�xq ~Osq ~w   ?@     q ~Axq ~�sq ~w   ?@     q ~�xq ~�sq ~w   ?@     q ~�q ~�q ~pxq ~sq ~w   ?@     q ~xq ~�sq ~w   ?@     q ~�xq ~$sq ~w   ?@     q ~Zq ~q ~^q ~ �xq ~�sq ~w   ?@     q ~�q ~yq ~0q ~�xq ~�sq ~w   ?@     q ~�xq ~wsq ~w   ?@     q ~jq ~Dxq ~ �sq ~w   ?@     q ~ �xq ~�sq ~w   ?@     q ~ �q ~�xq ~tsq ~w   ?@     q ~jxq ~ �sq ~w   ?@     q ~ �xq ~Ssq ~w   ?@     q ~Ixq ~sq ~w   ?@     q ~�q ~xq ~�sq ~w   ?@     q ~�xq ~�sq ~w   ?@     q ~�q ~xq ~�sq ~w   ?@     q ~wxq ~?sq ~w   ?@     q ~4q ~Uq ~�q ~�q ~�xq ~[sq ~w   ?@     q ~Qxq ~&sq ~w   ?@     q ~xq ~Fsq ~w   ?@     q ~<xq ~ �sq ~w   ?@     q ~ �xxsq ~ I?@     w      q ~ �sq ~w   @?@     q ~Hq ~�q ~:q ~hq ~�q ~�q ~(q ~�q ~ iq ~'q ~�q ~�q ~Dq ~ �q ~
q ~�q ~�q ~�q ~�q ~Aq ~�q ~zq ~�q ~�q ~jq ~$q ~�q ~Lq ~�xq ~ �sq ~w   @?@     #q ~ �q ~�q ~Qq ~�q ~q ~q ~�q ~\q ~"q ~�q ~yq ~q ~3q ~&q ~^q ~�q ~q ~�q ~�q ~q ~ �q ~ �q ~jq ~Iq ~q ~1q ~�q ~�q ~�q ~wq ~ �q ~q ~�q ~ �q ~xq ~7sq ~w   @?@     "q ~�q ~ Yq ~zq ~lq ~<q ~�q ~�q ~q ~ �q ~Uq ~Zq ~�q ~?q ~pq ~Nq ~�q ~ +q ~ �q ~fq ~�q ~�q ~pq ~q ~0q ~ qq ~]q ~�q ~�q ~ �q ~�q ~q ~/q ~�q ~�xq ~<sq ~w   ?@     q ~4q ~q ~ �q ~@q ~�q ~�q ~^q ~�q ~Vq ~zq ~�q ~�xxsq ~ I?@     w      q ~�sq ~w   ?@     q ~yq ~ q ~�q ~�xq ~nsq ~w   ?@     q ~iq ~2q ~�q ~�q ~q ~�xq ~�sq ~w   ?@     q ~�xq ~Usq ~w   ?@     q ~�q ~Pxxsr 5edu.cornell.cs.nlp.spf.base.hashvector.TreeHashVector�<�Lxs�� L valuest Ljava/util/TreeMap;xpsr java.util.TreeMap��>-%j� L 
comparatort Ljava/util/Comparator;xppw  �sq ~WD�t DYNSKIPppppsr java.lang.Double���J)k� D valuexr java.lang.Number������  xp��      sq ~W�"�q ~ t LEXt 0t 0psq ~n        sq ~W�"�q ~ q ~rt 0t 1psq ~n@$      sq ~W�&�q ~ q ~rt 1t 1psq ~n        sq ~W�މq ~ q ~rt 1t 10psq ~n@5oz�G�sq ~W�'qq ~ q ~rt 1t 7psq ~n@5oz�G�sq ~W�icq ~ q ~rt 10t 3psq ~n        sq ~W�i�q ~ q ~rt 10t 4psq ~n@$      sq ~Zw,hq ~ q ~rt 100t 11psq ~n�˃��>�sq ~Zvt�q ~ q ~rt 100t 5psq ~n?��H���sq ~Zvuq ~ q ~rt 100t 6psq ~n        sq ~ZvuPq ~ q ~rt 100t 8psq ~n�Ϣ�.��sq ~ZvxWq ~ q ~rt 101t 2psq ~n��.���.sq ~Zw3�q ~ q ~rt 102t 11psq ~n��8�8�sq ~Zw4	q ~ q ~rt 102t 12psq ~n        sq ~Zv|uq ~ q ~rt 102t 5psq ~n��xB�sq ~Zv�q ~ q ~rt 103t 0psq ~n?�J�a�sq ~Zv��q ~ q ~rt 104t 2psq ~n@�if�igsq ~Zv��q ~ q ~rt 105t 5psq ~n?�\��tsq ~Zv�q ~ q ~rt 105t 8psq ~n        sq ~Zv�q ~ q ~rt 106t 2psq ~n        sq ~Zv��q ~ q ~rt 107t 0psq ~n���5�#sq ~Zv�xq ~ q ~rt 107t 7psq ~n        sq ~Zv��q ~ q ~rt 108t 2psq ~n        sq ~Zv�_q ~ q ~rt 109t 2psq ~n        sq ~W�$�q ~ q ~rt 11t 12psq ~n        sq ~W�m�q ~ q ~rt 11t 6psq ~n@$      sq ~W�m�q ~ q ~rt 11t 8psq ~n        sq ~W�qaq ~ q ~rt 12t 7psq ~n@5oz�G�sq ~W�t�q ~ q ~rt 13t 3psq ~n@5oz�G�sq ~W�x)q ~ q ~rt 14t 1psq ~n@$      sq ~W�|Gq ~ q ~rt 15t 4psq ~n@$      sq ~W��q ~ q ~rt 16t 0psq ~n@$      sq ~W��q ~ q ~rt 16t 1psq ~n        sq ~Wă�q ~ q ~rt 17t 3psq ~n@5oz�G�sq ~Wă�q ~ q ~rt 17t 4psq ~n        sq ~WĈ%q ~ q ~rt 18t 9psq ~n@$      sq ~WĊ�q ~ q ~rt 19t 0psq ~n@,\��ў*sq ~WĊ�q ~ q ~rt 19t 1psq ~n@J�,��sq ~W�B�q ~ q ~rt 19t 10psq ~n�����z4sq ~Wċ�q ~ q ~rt 19t 7psq ~n�����sq ~W�*�q ~ q ~rt 2t 2psq ~n@5oz�G�sq ~W��eq ~ q ~rt 20t 0psq ~n�!pⴒ�sq ~W�݄q ~ q ~rt 20t 1psq ~n@:���h�qsq ~WŕVq ~ q ~rt 20t 10psq ~n�����|sq ~W��>q ~ q ~rt 20t 7psq ~n��@��)�sq ~W��q ~ q ~rt 21t 4psq ~n@$      sq ~WŜ�q ~ q ~rt 22t 11psq ~n@�F�ȑ�sq ~W��q ~ q ~rt 22t 5psq ~n@8r�t�u�sq ~W���q ~ q ~rt 22t 8psq ~n�!*�T�4Psq ~W��q ~ q ~rt 23t 3psq ~n@5oz�G�sq ~W��$q ~ q ~rt 23t 4psq ~n        sq ~W���q ~ q ~rt 24t 3psq ~n        sq ~W���q ~ q ~rt 24t 4psq ~n@$      sq ~W��q ~ q ~rt 25t 4psq ~n@$      sq ~Wū�q ~ q ~rt 26t 10psq ~n@5oz�G�sq ~W���q ~ q ~rt 26t 7psq ~n@5oz�G�sq ~W��	q ~ q ~rt 27t 3psq ~n@Al6sDsq ~W��(q ~ q ~rt 27t 4psq ~n@$      sq ~W���q ~ q ~rt 28t 2psq ~n@5oz�G�sq ~W��lq ~ q ~rt 29t 2psq ~n@5oz�G�sq ~W�.9q ~ q ~rt 3t 1psq ~n@$      sq ~W�Rq ~ q ~rt 30t 2psq ~n@5oz�G�sq ~W��q ~ q ~rt 31t 11psq ~n�!Q�8��sq ~W�V}q ~ q ~rt 31t 8psq ~n        sq ~W�Vq ~ q ~rt 32t 11psq ~n@xs��sq ~W�Y�q ~ q ~rt 32t 5psq ~n���Gf��sq ~W�Z>q ~ q ~rt 32t 8psq ~n@([@��٤sq ~W�Z]q ~ q ~rt 32t 9psq ~n        sq ~W�q ~ q ~rt 33t 11psq ~n?�W��#wsq ~W�]�q ~ q ~rt 33t 5psq ~n@��\?}sq ~W�]�q ~ q ~rt 33t 8psq ~n��Ɵ�sq ~W�`�q ~ q ~rt 34t 0psq ~n@E�/��sq ~W�`�q ~ q ~rt 34t 1psq ~n@/Q!u���sq ~W��q ~ q ~rt 34t 10psq ~n�!?�Ms�sq ~W�a�q ~ q ~rt 34t 7psq ~n@ �^n��sq ~W��q ~ q ~rt 35t 11psq ~n@�+;�Y,sq ~W�eCq ~ q ~rt 35t 6psq ~n        sq ~W� Zq ~ q ~rt 36t 11psq ~n@ ����sq ~W�h�q ~ q ~rt 36t 5psq ~n        sq ~W�iBq ~ q ~rt 36t 8psq ~n�&���sq ~W�lIq ~ q ~rt 37t 2psq ~n��,�\2��sq ~W�p
q ~ q ~rt 38t 2psq ~n?�o�r9�sq ~W�s�q ~ q ~rt 39t 2psq ~n@/4g��sq ~W�28q ~ q ~rt 4t 3psq ~n@5oz�G�sq ~W��aq ~ q ~rt 40t 2psq ~n���=J�sq ~W��"q ~ q ~rt 41t 2psq ~n@"9!rsq ~W���q ~ q ~rt 42t 2psq ~n�+L0�0�sq ~W��fq ~ q ~rt 43t 0psq ~n@�X�Xsq ~W�хq ~ q ~rt 43t 1psq ~n��,��,�sq ~W��'q ~ q ~rt 44t 0psq ~n�8��8��sq ~W��Fq ~ q ~rt 44t 1psq ~n@r�*r�*sq ~Wƍq ~ q ~rt 44t 10psq ~n        sq ~W���q ~ q ~rt 45t 0psq ~n        sq ~W���q ~ q ~rt 46t 2psq ~n@.ffffffsq ~WƘzq ~ q ~rt 47t 11psq ~n���o��sq ~W��bq ~ q ~rt 47t 8psq ~n@.ffffffsq ~W��q ~ q ~rt 47t 9psq ~n        sq ~W��+q ~ q ~rt 48t 0psq ~n?����t�sq ~W��Jq ~ q ~rt 48t 1psq ~n        sq ~WƜq ~ q ~rt 48t 10psq ~n���,�3�sq ~W��q ~ q ~rt 48t 7psq ~n��(C�Isq ~WƟ�q ~ q ~rt 49t 11psq ~n������sq ~W��q ~ q ~rt 49t 9psq ~n        sq ~W�5�q ~ q ~rt 5t 2psq ~n@5oz�G�sq ~W�;q ~ q ~rt 50t 5psq ~n��YL�sq ~W�;zq ~ q ~rt 50t 8psq ~n@ �LE�jsq ~W�;�q ~ q ~rt 50t 9psq ~n        sq ~W�>Cq ~ q ~rt 51t 0psq ~n@rPt^�sq ~W�>bq ~ q ~rt 51t 1psq ~n��ŕ��sq ~W��4q ~ q ~rt 51t 10psq ~n��e���sq ~W�?q ~ q ~rt 51t 7psq ~n��o�sq ~W�Bq ~ q ~rt 52t 0psq ~n@�I+}G�sq ~W�B#q ~ q ~rt 52t 1psq ~n��9�Be�isq ~W���q ~ q ~rt 52t 10psq ~n���'?b:�sq ~W�B�q ~ q ~rt 52t 7psq ~n@ٳN�Dsq ~W�Fq ~ q ~rt 53t 2psq ~n@t!	�sq ~W�I�q ~ q ~rt 54t 2psq ~n?���l��sq ~W�MGq ~ q ~rt 55t 0psq ~n@$��c��sq ~W�Mfq ~ q ~rt 55t 1psq ~n����;5Y)sq ~W�8q ~ q ~rt 55t 10psq ~n�vEҦBsq ~W�N q ~ q ~rt 55t 7psq ~n�"�Au���sq ~W�QFq ~ q ~rt 56t 2psq ~n@       sq ~W�Uq ~ q ~rt 57t 2psq ~n�l8���2sq ~W�X�q ~ q ~rt 58t 0psq ~n�,�)S�
sq ~W�X�q ~ q ~rt 58t 1psq ~n���fxܪsq ~W�{q ~ q ~rt 58t 10psq ~n�)I�gesq ~W�Ycq ~ q ~rt 58t 7psq ~n@7����sq ~W�\�q ~ q ~rt 59t 2psq ~n        sq ~W�9�q ~ q ~rt 6t 3psq ~n@5oz�G�sq ~W�gq ~ q ~rt 60t 12psq ~n        sq ~WƳ=q ~ q ~rt 61t 5psq ~n        sq ~Wƶ�q ~ q ~rt 62t 2psq ~n@f�}�Ogsq ~W�r4q ~ q ~rt 63t 11psq ~n�.ffffffsq ~W�rSq ~ q ~rt 63t 12psq ~n        sq ~Wƾ#q ~ q ~rt 64t 2psq ~n�2�Γ*�sq ~W���q ~ q ~rt 65t 2psq ~n?�� ��FHsq ~W��!q ~ q ~rt 66t 6psq ~n        sq ~W��fq ~ q ~rt 67t 2psq ~n��#"5��sq ~WǄ�q ~ q ~rt 68t 11psq ~n?�.���*sq ~W�̈́q ~ q ~rt 68t 5psq ~n        sq ~W���q ~ q ~rt 69t 2psq ~n@�}�{ lsq ~W�=q ~ q ~rt 7t 0psq ~n@$      sq ~W�==q ~ q ~rt 7t 1psq ~n        sq ~W��Pq ~ q ~rt 70t 11psq ~n?�      sq ~W��oq ~ q ~rt 70t 12psq ~n        sq ~W�#�q ~ q ~rt 70t 5psq ~n�       sq ~W�$8q ~ q ~rt 70t 8psq ~n?�      sq ~W��q ~ q ~rt 71t 11psq ~n?�      sq ~W�'�q ~ q ~rt 71t 5psq ~n��      sq ~W�(q ~ q ~rt 71t 9psq ~n        sq ~W�+ q ~ q ~rt 72t 2psq ~n        sq ~W�.�q ~ q ~rt 73t 0psq ~n@�9�P��sq ~W�.�q ~ q ~rt 73t 1psq ~n�-��l��nsq ~W��tq ~ q ~rt 73t 10psq ~n��      sq ~W�/\q ~ q ~rt 73t 7psq ~n��T4��sq ~W��Tq ~ q ~rt 74t 11psq ~n?�6?�'�sq ~W�2�q ~ q ~rt 74t 5psq ~n��.���.sq ~W�2�q ~ q ~rt 74t 6psq ~n        sq ~W�3<q ~ q ~rt 74t 8psq ~n@�8�;sq ~W�7q ~ q ~rt 75t 9psq ~n        sq ~W�:�q ~ q ~rt 76t 6psq ~n        sq ~W�>Aq ~ q ~rt 77t 6psq ~n        sq ~W�A�q ~ q ~rt 78t 2psq ~n��������sq ~W��8q ~ q ~rt 79t 12psq ~n        sq ~W�A[q ~ q ~rt 8t 4psq ~n@5oz�G�sq ~WǗ�q ~ q ~rt 80t 2psq ~n�0�'U��sq ~Wǜq ~ q ~rt 81t 6psq ~n        sq ~Wǟ!q ~ q ~rt 82t 0psq ~n��x�y�;sq ~Wǟ@q ~ q ~rt 82t 1psq ~n        sq ~Wǣ q ~ q ~rt 83t 2psq ~n?��Q��sq ~W�^�q ~ q ~rt 84t 11psq ~n��Πq��sq ~Wǧ�q ~ q ~rt 84t 8psq ~n�!�|�=�sq ~WǪ�q ~ q ~rt 85t 2psq ~n@�_2�G�sq ~WǮ%q ~ q ~rt 86t 0psq ~n?��f��sq ~WǮDq ~ q ~rt 86t 1psq ~n        sq ~Wǲ�q ~ q ~rt 87t 5psq ~n��      sq ~Wǲ�q ~ q ~rt 87t 6psq ~n        sq ~Wǲ�q ~ q ~rt 87t 8psq ~n��      sq ~Wǵ�q ~ q ~rt 88t 0psq ~n����h��sq ~W�m�q ~ q ~rt 88t 10psq ~n        sq ~WǶ�q ~ q ~rt 88t 7psq ~n��8�8�sq ~Wǹhq ~ q ~rt 89t 0psq ~n��8�8�sq ~Wǹ�q ~ q ~rt 89t 1psq ~n�,O�E�]sq ~W�qYq ~ q ~rt 89t 10psq ~n��;�jSsq ~WǺAq ~ q ~rt 89t 7psq ~n��8�Fz�2sq ~W���q ~ q ~rt 9t 11psq ~n@5oz�G�sq ~W���q ~ q ~rt 9t 12psq ~n@5oz�G�sq ~W�E;q ~ q ~rt 9t 5psq ~n        sq ~W��q ~ q ~rt 90t 0psq ~n���
�ѧrsq ~W�q ~ q ~rt 90t 1psq ~n        sq ~W��q ~ q ~rt 90t 7psq ~n��!0�V�sq ~W��q ~ q ~rt 91t 2psq ~n?�������sq ~W��q ~ q ~rt 92t 2psq ~n@ �oq��psq ~W��Qq ~ q ~rt 93t 11psq ~n���g�sq ~W��q ~ q ~rt 93t 5psq ~n        sq ~W�9q ~ q ~rt 93t 8psq ~n?��g�sq ~W��q ~ q ~rt 94t 11psq ~n���f����sq ~W��q ~ q ~rt 94t 5psq ~n?��f����sq ~W�q ~ q ~rt 94t 9psq ~n        sq ~W���q ~ q ~rt 95t 11psq ~n���f����sq ~W���q ~ q ~rt 95t 12psq ~n        sq ~W�^q ~ q ~rt 95t 5psq ~n?��f����sq ~W�ڔq ~ q ~rt 96t 11psq ~n���f����sq ~W�#q ~ q ~rt 96t 5psq ~n?��f����sq ~W�#>q ~ q ~rt 96t 6psq ~n        sq ~W�&Eq ~ q ~rt 97t 0psq ~n        sq ~W�&dq ~ q ~rt 97t 1psq ~n?�/p&��.sq ~W��6q ~ q ~rt 97t 10psq ~n��bv'bv'sq ~W�'q ~ q ~rt 97t 7psq ~n@��r�sq ~W�*%q ~ q ~rt 98t 1psq ~n��y�԰asq ~W���q ~ q ~rt 98t 10psq ~n���;�;sq ~W�*�q ~ q ~rt 98t 7psq ~n�	#0#0sq ~W�.bq ~ q ~rt 99t 5psq ~n?�y~�?*sq ~W�.�q ~ q ~rt 99t 6psq ~n@1c1cq ~sq ~n?�      sq ~e��q ~ t TMPt 0ppsq ~n?��H�ӝ�sq ~e���q ~ q ~
�t 1ppsq ~n        sq ~e�A>q ~ q ~
�t 10ppsq ~n�}!���sq ~e�D�q ~ q ~
�t 11ppsq ~n��Z[F�fVsq ~e�H�q ~ q ~
�t 12ppsq ~n        sq ~e��q ~ q ~
�t 2ppsq ~n?�16	V�sq ~e�Rq ~ q ~
�t 3ppsq ~n?�AC�W�sq ~e�
q ~ q ~
�t 4ppsq ~n        sq ~e��q ~ q ~
�t 5ppsq ~n?�^V�EJ�sq ~e��q ~ q ~
�t 6ppsq ~n?�x'�x'�sq ~e�Vq ~ q ~
�t 7ppsq ~n?�c�8ɀ�sq ~e�q ~ q ~
�t 8ppsq ~n        sq ~e��q ~ q ~
�t 9ppsq ~n        q ~sq ~n?�      sq ~{H�q ~ t XEMEt 0ppsq ~n@$      sq ~{H��q ~ q ~
�t 1ppsq ~n@$      sq ~{^�0q ~ q ~
�t 10ppsq ~n@$      sq ~~��q ~ q ~
�t 100ppsq ~n?�+R5�Lsq ~~�Cq ~ q ~
�t 101ppsq ~n��.���.sq ~~q ~ q ~
�t 102ppsq ~n���[�!�sq ~~�q ~ q ~
�t 103ppsq ~n?�J�a�sq ~~�q ~ q ~
�t 104ppsq ~n@�if�igsq ~~Gq ~ q ~
�t 105ppsq ~n?�\��tsq ~~q ~ q ~
�t 106ppsq ~n        sq ~~�q ~ q ~
�t 107ppsq ~n���5�#sq ~~�q ~ q ~
�t 108ppsq ~n        sq ~~Kq ~ q ~
�t 109ppsq ~n        sq ~{^��q ~ q ~
�t 11ppsq ~n@$      sq ~{^��q ~ q ~
�t 12ppsq ~n@$      sq ~{^�sq ~ q ~
�t 13ppsq ~n@$      sq ~{^�4q ~ q ~
�t 14ppsq ~n@$      sq ~{_ �q ~ q ~
�t 15ppsq ~n@$      sq ~{_�q ~ q ~
�t 16ppsq ~n@$      sq ~{_wq ~ q ~
�t 17ppsq ~n@$      sq ~{_8q ~ q ~
�t 18ppsq ~n@$      sq ~{_�q ~ q ~
�t 19ppsq ~n@$      sq ~{H��q ~ q ~
�t 2ppsq ~n@$      sq ~{_b�q ~ q ~
�t 20ppsq ~n@,綛f7|sq ~{_fPq ~ q ~
�t 21ppsq ~n@$      sq ~{_jq ~ q ~
�t 22ppsq ~n@$      sq ~{_m�q ~ q ~
�t 23ppsq ~n@$      sq ~{_q�q ~ q ~
�t 24ppsq ~n@$      sq ~{_uTq ~ q ~
�t 25ppsq ~n@$      sq ~{_yq ~ q ~
�t 26ppsq ~n@$      sq ~{_|�q ~ q ~
�t 27ppsq ~n@. ��9�sq ~{_��q ~ q ~
�t 28ppsq ~n@$      sq ~{_�Xq ~ q ~
�t 29ppsq ~n@$      sq ~{H�Dq ~ q ~
�t 3ppsq ~n@$      sq ~{_��q ~ q ~
�t 30ppsq ~n@$      sq ~{_گq ~ q ~
�t 31ppsq ~n�!Q�8��sq ~{_�pq ~ q ~
�t 32ppsq ~n@,1�]y�rsq ~{_�1q ~ q ~
�t 33ppsq ~n��pjD�sq ~{_��q ~ q ~
�t 34ppsq ~n@2�sozsq ~{_�q ~ q ~
�t 35ppsq ~n@�+;�Y,sq ~{_�tq ~ q ~
�t 36ppsq ~n���g�";sq ~{_�5q ~ q ~
�t 37ppsq ~n��,�\2��sq ~{_��q ~ q ~
�t 38ppsq ~n?�o�r9�sq ~{_��q ~ q ~
�t 39ppsq ~n@/4g��sq ~{H�q ~ q ~
�t 4ppsq ~n@$      sq ~{`KMq ~ q ~
�t 40ppsq ~n���=J�sq ~{`Oq ~ q ~
�t 41ppsq ~n@"9!rsq ~{`R�q ~ q ~
�t 42ppsq ~n�+L0�0�sq ~{`V�q ~ q ~
�t 43ppsq ~n��Y��Y��sq ~{`ZQq ~ q ~
�t 44ppsq ~n?�Y��Y��sq ~{`^q ~ q ~
�t 45ppsq ~n        sq ~{`a�q ~ q ~
�t 46ppsq ~n@.ffffffsq ~{`e�q ~ q ~
�t 47ppsq ~n@)8�J�e�sq ~{`iUq ~ q ~
�t 48ppsq ~n�!�\����sq ~{`mq ~ q ~
�t 49ppsq ~n������sq ~{H��q ~ q ~
�t 5ppsq ~n@$      sq ~{`��q ~ q ~
�t 50ppsq ~n@
�~���sq ~{`�mq ~ q ~
�t 51ppsq ~n����%|(�sq ~{`�.q ~ q ~
�t 52ppsq ~n@�j����sq ~{`��q ~ q ~
�t 53ppsq ~n@t!	�sq ~{`ΰq ~ q ~
�t 54ppsq ~n?���l��sq ~{`�qq ~ q ~
�t 55ppsq ~n�"h{8��sq ~{`�2q ~ q ~
�t 56ppsq ~n@       sq ~{`��q ~ q ~
�t 57ppsq ~n�l8���2sq ~{`ݴq ~ q ~
�t 58ppsq ~n@�h#�`sq ~{`�uq ~ q ~
�t 59ppsq ~n        sq ~{H��q ~ q ~
�t 6ppsq ~n@$      sq ~{a4q ~ q ~
�t 60ppsq ~n        sq ~{a7�q ~ q ~
�t 61ppsq ~n        sq ~{a;�q ~ q ~
�t 62ppsq ~n@f�}�Ogsq ~{a?Nq ~ q ~
�t 63ppsq ~n�.ffffffsq ~{aCq ~ q ~
�t 64ppsq ~n�2�Γ*�sq ~{aF�q ~ q ~
�t 65ppsq ~n?�� ��FHsq ~{aJ�q ~ q ~
�t 66ppsq ~n        sq ~{aNRq ~ q ~
�t 67ppsq ~n��#"5��sq ~{aRq ~ q ~
�t 68ppsq ~n?�.���*sq ~{aU�q ~ q ~
�t 69ppsq ~n@�}�{ lsq ~{H�Hq ~ q ~
�t 7ppsq ~n@$      sq ~{a�jq ~ q ~
�t 70ppsq ~n        sq ~{a�+q ~ q ~
�t 71ppsq ~n        sq ~{a��q ~ q ~
�t 72ppsq ~n        sq ~{a��q ~ q ~
�t 73ppsq ~n� ݲ$��sq ~{a�nq ~ q ~
�t 74ppsq ~n@�n��sq ~{a�/q ~ q ~
�t 75ppsq ~n        sq ~{a��q ~ q ~
�t 76ppsq ~n        sq ~{a±q ~ q ~
�t 77ppsq ~n        sq ~{a�rq ~ q ~
�t 78ppsq ~n��������sq ~{a�3q ~ q ~
�t 79ppsq ~n        sq ~{H�	q ~ q ~
�t 8ppsq ~n@$      sq ~{b�q ~ q ~
�t 80ppsq ~n�0�'U��sq ~{b �q ~ q ~
�t 81ppsq ~n        sq ~{b$Kq ~ q ~
�t 82ppsq ~n��x�y�;sq ~{b(q ~ q ~
�t 83ppsq ~n?��Q��sq ~{b+�q ~ q ~
�t 84ppsq ~n�"�f����sq ~{b/�q ~ q ~
�t 85ppsq ~n@�_2�G�sq ~{b3Oq ~ q ~
�t 86ppsq ~n?��f��sq ~{b7q ~ q ~
�t 87ppsq ~n�       sq ~{b:�q ~ q ~
�t 88ppsq ~n� צq¢�sq ~{b>�q ~ q ~
�t 89ppsq ~n�2�sozsq ~{H��q ~ q ~
�t 9ppsq ~n@$      sq ~{b�(q ~ q ~
�t 90ppsq ~n��n��(R�sq ~{b��q ~ q ~
�t 91ppsq ~n?�������sq ~{b��q ~ q ~
�t 92ppsq ~n@ �oq��psq ~{b�kq ~ q ~
�t 93ppsq ~n        sq ~{b�,q ~ q ~
�t 94ppsq ~n        sq ~{b��q ~ q ~
�t 95ppsq ~n        sq ~{b��q ~ q ~
�t 96ppsq ~n        sq ~{b�oq ~ q ~
�t 97ppsq ~n@P�9:�sq ~{b�0q ~ q ~
�t 98ppsq ~n�P�9:�sq ~{b��q ~ q ~
�t 99ppsq ~n@��"mP�q ~sq ~n?�      sq ~��.�t LOGCOOCt ARGARGq ~ �q ~ �psq ~n?Φ�$��sq ~�ȃq ~Aq ~Bq ~�q ~ �psq ~n�%�M�ـTsq ~�l*�q ~Aq ~Bq ~�q ~�psq ~n���k��sq ~�$��q ~Aq ~Bq ~ Bq ~ �psq ~n@"�9���#sq ~��9fq ~Aq ~Bq ~ Bq ~�psq ~n��9��Jsq ~�>΃q ~Aq ~Bq ~ Bq ~ Bpsq ~n��vm�xvsq ~�>��q ~Aq ~Bq ~qq ~ �psq ~n@=�N阤sq ~�↨q ~Aq ~Bq ~qq ~�psq ~n�%��QhPsq ~�Y�q ~Aq ~Bq ~qq ~ Bpsq ~n@dە nsq ~J�Cq ~Aq ~Bq ~qq ~qpsq ~n� ����sq ~N�q ~Aq ~Bq ~�q ~ �psq ~n�/�?'K�sq ~�d�q ~Aq ~Bq ~�q ~�psq ~n����>��sq ~h�q ~Aq ~Bq ~�q ~ Bpsq ~n���8*isq ~����q ~Aq ~Bq ~�q ~qpsq ~n?���>���sq ~�E-q ~Aq ~Bq ~�q ~�psq ~n@#��L�Nsq ~�
��q ~Aq ~Bt varq ~�psq ~n�!M�9��sq ~�q ~At PREDARGq ~ Eq ~apsq ~n@W����sq ~vF8uq ~Aq ~dq ~�q ~ �psq ~n@"a�=Musq ~+��Vq ~Aq ~dq ~�q ~�psq ~n�-��W���sq ~�`usq ~Aq ~dq ~�q ~ Bpsq ~n@$w`j.sq ~�w�q ~Aq ~dq ~�q ~qpsq ~n?�Jm���sq ~Ę�gq ~Aq ~dq ~�q ~�psq ~n?�1u{��sq ~Epf'q ~Aq ~dq ~ �q ~apsq ~n����2W�sq ~$�"Bq ~Aq ~dq ~�q ~�psq ~n�>�-VϚsq ~DA�fq ~Aq ~dq ~�q ~apsq ~n�-��W���sq ~0"0�q ~Aq ~dq ~ Bq ~�psq ~n@*�7��3�sq ~O���q ~Aq ~dq ~ Bq ~apsq ~n@$w`j.sq ~Q�+q ~Aq ~dq ~qq ~apsq ~n�#��e�sq ~q��q ~Aq ~dq ~ xq ~�psq ~n@I�>�\fsq ~�k�uq ~Aq ~dq ~�q ~apsq ~n�$��4Lsq ~���q ~Aq ~dq ~�q ~ Epsq ~n@W����sq ~T�ڒq ~Aq ~dq ~�q ~�psq ~n���8���sq ~(�yq ~Aq ~dq ~�q ~ �psq ~n��(j��lsq ~��@�q ~Aq ~dq ~�q ~qpsq ~n�>2k��C�sq ~w!qkq ~Aq ~dq ~�q ~�psq ~n�,�cV���sq ~k#�t LOGEXPt CPAPq ~�q ~�t 1sq ~n��UUUUUUsq ~Β��q ~�q ~�q ~�q ~ Bt 1sq ~n�"/��4�msq ~���q ~�t CPP1q ~�q ~ Bq ~�sq ~n�������sq ~(��-q ~�q ~�q ~�q ~qq ~ �sq ~n@=�N阤sq ~�Σq ~�q ~�q ~�q ~�q ~ �sq ~n�/�?'K�sq ~D��q ~�q ~�q ~�q ~�q ~qsq ~n?���>���sq ~�רq ~�t REPTq ~�q ~ �psq ~n?Φ�$��sq ~r��q ~�q ~�q ~�q ~�psq ~n��B�Y!dsq ~� �q ~�q ~�q ~�q ~ Bpsq ~n@ٳN�Dsq ~(�$q ~�q ~�q ~�q ~qpsq ~n� ����sq ~XG�q ~�q ~�q ~�q ~�psq ~n@#��L�Nsq ~d!+�t RULEt <applypppsq ~n?�1c1csq ~��	�q ~�t >applypppsq ~n@#gT~�sq ~"A�q ~�t >comp1pppsq ~n��35���sq ~4::�q ~�t 	>thatlesspppsq ~n�#-����x